`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
KPwPdORyW3jQITxLU49ITpHIAc2EUwMUYAoRqiVUfUeZHTBvElxtzMD0AHIkDItAix/LyOCXDC1z
lGVPLedIHQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
gsUAYdj8+YC1BLMqJksFvsSUcBCneybpvDdqbaHRbG1FQ64ag+QXCA3uwhj35S0PY71NGGygS5ur
7QAVZae0Qx1cxiaGQMN1Y1VbvrH/EBsPdjpyzc8LwZKUkvDTZi4KDPT/sqrfucrYavLnzIjv695n
FMoh8a+9jn3QAgoEwD8=

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
q+XzY0hwi2oRHlU9ipRQM5109658PZKlTdYyF2I4rYki5o3rP2AgHHK+2FWeyRkBz2Pi3MvOjmeH
Puez3oeZA5OMacY0fn0hVEb2A7gFZc8m2y/5pZ430MlzJ+c63yC3bARPK/djDr+BaK6q2OtiNAaC
Edh9rtN/YRfvDOT8ElM=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
D1bwrBkg1d9MGz/3Bx6L9m8zNqWzXs7en1acM4DcH7Ig2bZX+ZU8qanwUDwYG+uQqPPU/eTX4Anv
ffcg4mYQgmUDQVAmtWpU5dyuq1HgaXelTWY9nvFSQHDKSz8H1FhFOXa+J68fYXQyABgULkdfW6Nv
SQIilL16bUH9ue+BB8D4tNTYkJ/jq6z9/F10H75raT0S7nWksRzFk1N/5zYtcXIgsLhajVmVyxAg
y9J6tPkHSs68iw5AQcqxQ/HzuMhC6d+TXwe6v6teitp3BPxZxBd68GOOJ1ZKkmuEvoqHkjghy3yx
LJXqNBjX6toptbVvJTBynH9qSWBlYv3t6NO7/Q==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
k2YBUjEJGyp0+OR5dN1t6doID6L1rLo44M1w0g1RmPKAToarp+Y83ga1s+j+Gkv/eF0m9JIYhtXU
mhOB5v5djBfAMQ39h65dDVtmTtqq3OW5HSOHN9rMcqStpV927AS+hftD8zwu9BZbERxpKc29KiQz
81pBJALmXJoiVKoUvaawzO+bfgNm+E9dZnaX5G5NKLWSxfMrJwLzkVyCEmBT+Jm3s0Jwe9pD8Rjr
lbEg/GugQytMJ7X75dVQlleUwA3IruTPBng8hC62+C5eb5fbargQ9D4wyuDXTQMIS79uxk1f/6e7
yv5Fntv24HgV8zZ/PRzP4KackR+Mjpz8oB8mGQ==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
IOjxX1MzevlKWK3S2QEhgC0hId6CVQ+BtQPo8WqeBkCu94/1dpI08VQKsCaqY1NIDXE6S5vvmHRU
JqpFAwdQeBt5zpD68kvsDgwM/HNFVyzqaAm/QI9lEfPhUEBOuLdu0hva6MTXFgt9agFfQIsC+a0J
YmxxlzlJ3LB0wl+n4r1N/3naMofMSEx48vxBdbzdOqhUFwUaQ4TWqTzKfVsJLp3WiI7nBAvz4Fbj
5MjA+QPRFWcj9BKy8VqFQk9+f0iUZ1x9qmjk8AL5+QxkFVT4WjwDNk3zSUgvqH0dM7Bi8lHSHNqS
miFEFHstFHTJF3MPalhgTojxpWiJeqnXp/zPvQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 779648)
`protect data_block
7MIbn+VTupd25XoYfTNSEco+iVs/4DQmxN/3cDxiwH4X0GnEaqT3Nj3it28x/VFDg80dr52lWylR
JV7F/mY0F7vN/hYAaPr4Q4gOSO6ZFn9AEOQwmhGaQSyk9Dguj++HLOT0BVtiwL4vlD1hL1dS7HBW
bRcQWBxuYUpO++6eysUaDyeJ1H/1SMZwpr8Oy14EG6GorZ069RRgGPjsrKbVGZM53WToReB5pd3c
IyeUzn9yWoZNgmMY7zo3kzDjyp22FU5zcn5yVd8D+eA4SEV6RuqdhGhKtUKDq76/fKjObL4RX4zx
nDWl8rgcDNUNmaigFkWiv07wFxqe8YcC7WaGM9AI3dJwfmMZzZ4ZqhqXbAHJ+hiCFWhAuMe9DRqI
jtIE/mUQ/olI55vNpAVKG7ZO1CH9yaydos76Fgy9/2aoN8YLap+efseaOL+tRgu3t1LMU2gfHbzJ
0DbbbTNhD5/IOEzoWn5F+0KAfEDsCi8slWe+xBmVxley4INct2x1DXdwDL6CH6UzEUqyI9mEthUa
tQcCuh6miaECjlzb0oPLNBfEL1CDLN43HDPLpjTxTO5N1gurN67vcgapcWNhn735I+jYebblLP36
4VsH4F6qwAWGbHIaIqx4vFhLhjWYTUGCqT12ePrcGZ44dai/vzjRGOFdU8y7pUz0XMQ2xa9lW949
9qlv9wePItppG+SCYYRr5usPsSq+NfH1n2cKUwsszDhc0XN53ekNQaj9rOnO37+P2JSFqCblZgL/
9O4tw3IR2x6r7ROSsyh9Gitm5ED86AGhIybGe6OR0ABdZawwO8/0rLpbI8VLY9hFjg2WpOlCENvL
AB09qi05Tc3G9t60Qajq2HmhSy2XWvtU3/QePHvH7CtopEFCBENsXGy4dyjBf+XisjRS3QQEEQSB
0sG3tcyXJfoQkPgUqt7XSzbZJ8lvh8r61TE4nLE7LfUyZT5fxIvu2XkkedgkvzxXyqcYVueLG9Rm
YF3xLYe4RDmY6r2UvUzz+Mjkv7zQSMDwbWJKQ1z9v5MK+gLbt+1bgUQetO2gfr0kHcDrr0stQMux
qKuDOfq12VowLQrheqoD1OlDtef5uBU6EcxjIPX7adK4RTY1n8ohxWV7S6gUZSlWMrOT/cPNFNce
UV2toTDedjoNWOfJOq2WlsB8H6ZOGFKHBOgG6gdEbd6C/BLgVeWl3Z7sDt3eLAsP5lVAb6trgdZc
pwu18TRD/V/UkevXOpTLJDCTqLvSwgPV1h7Ls9OJzuOXx/IJHXtVFpTx7RO0afu2K96MRpRL3eoU
2sfG4WOA0dlThp5uykx5t0hHAnojXJ3kEIlDEoStvQ9tmr6oDhjUjrKHAQ0E4T/baaPlRZN5xZMg
tI2wgMiSJVWW/V0bnGK0lFTzcVJQkorjY3ScY752w474HY/9CPcaP1yZUWYivls6fT+Sirjt20di
IvQ7VMWCrOVLpM1Hz1mkgJkfTv59yjKUB0YhvxJnERmpZyOKcolvxl3OA8WnpjHQcrrPqbU2U4FD
Od1X4QsL09WA+y/tfFJt6fsunS1fVHI3GrzsmDXwA/KnafUXJT/EzdMHMXNNUiSKW/Bh/zHOLQbq
BYxL+3fNsjcKArZ7R6JK3vQD5AJzqEXMjBws/LaMIr4lQiZOQ6W3zxuGot+sdfmmF+HJVXxbwqAX
OId10/iR834oAQ5aEJYXXgiy9IDVPFPjxvD2c3dtGce3TSu5aQISGDpm9O9YFER6BzcXe5CJ2qrp
EsQLgCP2IHGqB0ekN7NGFp2HYTnoaL4CMa6fpbpFaJrgW/0LlRBILJUEoKxNlVEmTf/QArze594r
N/BzZEi1lQVQzAkQR/UPPzPpiuODq/lgCtInZD55AMwCU/DP76fWA6o7vVTWe1xFnvq1l6E+Jml/
W+YnO0Z9J+0yDpGAjWOCiJhJomzvVqDNqk94x8flfafYY5W4ZHuoekbX8Szd8aUr6V+S+lr+Ma+J
a/eUw7cVhyfQISv0lKYzFjAks0+1Wp0G8Jx5RFZsBMmxDjXBuDIZ5KJip1QM4qggJ9fcZa7hKulN
QLKwOnOseMGmq9lzXBA8QG3Q/k+iGwRBZIJyilKKXKW38LiC/ZyyYG0sbgXKDJWU+U4dhUw2F+Zc
8EpMhXXOTWHGByoZjttH32Oq5OBqyyEpzDH1ETrU/q2Q3QsSkQyyOnm/uMIHL9MB5k2NgqyQXN3v
tx/JOXFk5eP+vQ/lUW3MJ8bRjPpcmhuOn/m3hJrU/aNZlvgSxpuexoIotHc4VZLISF8hqVTcQo+V
YEcHDxISZ7FmXaix+Bk/VFOeyfCGanfRIZh2P+6wPpxnVkOn78P0SAieg5DzuDBHZFRClpYnGYdH
v6lOeLRLAKJJUpO1MqK6Q/O+2BFGBK4f7MFIgH9zy1clrhbZmnH7US6AwMa9lu+uxnXPNvGEaL1V
IRRLuNDDBtf2SVNps6YiBmOimYWWLTIIF4LnNL8szO7y1YsLd79YOZncN7/sxrIj+VBFpdkhR38h
BpjFbKOjJyeIV2YO3DzBSBp/3espgKNwUv9sDThdD7lQZ7a2lptns6G2bCocAzZKydJO6iOm4mfa
GAfxgClzH1XKEo7t31u54CRJj9CW1X0ntScjapi0hVZQonJt3W98cUuXhBlhRLg7I1vlqZvQKsZQ
+UGIklmwz+c4yzuRX7CcEG+Vo3p5RRvgCLhRm7apg86iY2eW7uzNdaRk0monxf/qDlWCLlfznTiE
v+DY7YNGo8pAY+UEpYcGI2WheKTylHdqtjSISZZVOC49eOnlSTdK9pP38nUOeVW95BCOJ8cNwKDd
h+mq4NsQzJTpDFUquOAJenSBR3vvmJTUwPn58DoMSKBo8A3kwDPlL7oKFkZn81IA1fvl8+8NLDRY
9dJOjpDuzmdbQiHoYiPecBLJYM3owaYNr97DBYaUC6VS6MJ9swJFPKOpltmNWSRgv1eI/7W2MPNc
uw+k3diMPiEWNM3PjkWS1vDmqmMq7CW25f8/4Z+JORDVJu+f9tJUMnQm4gq76rwo6HS4llLh1sHQ
zDcfY41rrZMX4yyM0QUWFdJUtynVMyXAoWzGxOS86lSwJXgRUUqBAw7JGDzxY1xv4AItAinMChj3
iAZ6gquN9sh42y48rSMYeLcCLYClTKTWmoH/aIFtcYRBv520cPOv/0zz0uIQXyx8UPGv+xrF7Y9q
/5f1yteonwqZ9rvWgj9BbA6Q4cZuCy/D6fy3K0M1X4dOdcxGhl1qVHhMcy5I6LUcUeX1UIhSmtYK
k8t0/KIa5zL4MPvBIZjhHAs4E+6q/sEs0Ev27jGl9JKeN56uwsy8yJkIKh3V1TrSJsqow65otZcD
0rVo9uK7bhI0uEyat0dcuOYy2ipqm6LFRxR25MjaQnW+PBPYZWxrjStELsKDWVLH3J3OWlfDu+FQ
nQ7mOXeaw4Am04//yDxp+ab9q5crEPpHHKPoNCMHmUX9o5z3tB05E8g+3ER7qFIWb5fbYiZ9elwb
n1VVrBHAmVSqd6uv9Fy0tMsTqV8nLdOL5j0uR39MjduXZTZZWpTbm6gDcdqjrnDkM+ucvQyx8ZhO
cm75gfbnRUdGma6ciXHMX2IHhChDKV4rdiGoudcA6ZMjD4YroqCeborTUyuE4ncIdj0OJXstWjAB
JiKaechnS1OeFKa0OFE0gOUYjGAb97zjljvvPWc+WFK7XLhABEvYnsIC4CMIx8u6nyVc0s7WZOKL
XoPDWnGSYU94OVY/wAaqDT7aJw7oqUgMIIU9CcrOsrCkbKdJGV5vgtFOZTO3Yp7wuVEHhtLBB/+t
c7nHNM6xDeN604GJ0K/7MjiSrcq08/il+Ta9O2GKajUTpKclE3EdLmStQdxZ457sb0qpjulEbZIl
8u2Ah8KkWyY589wXf1fMHjv9Pz+78HMkSQiRGCCcg16XXsxB4DoRfBmHVMMgaAK6O6ADrdTl2QSv
ndojoVJsO9Yeeexv5ZxNleJj1V6g/OWUVQV5JZll6w87S43F6NuMW0eWYxTxuI2g2t692akzi7WY
lTxqNNUUQNQngzIIIui3NJ5Ahw0kVh4IbCqS/L/VNEHA3zjTA/ZiWxe2a9B/r/pJChPIxynFB4xa
mlt9SF51ktRoagVkCvl6lVf6/KyoUCQRWAaWzM6WxN6b4kFZd7m4XT727tKrAiuIf9oWx0Dllkn3
rBLdYt9yriGY2g+ciw/hIOzJ1T2hzkuXG73nlK5pf5Dnlcy1RKapsgHWN29wcrg3K+zdgZ6JSMAr
IyQSYryXBmWARzRw5FJlydMUQd87xt/IgGOjVb/eZFXp4pd3n6wZ/sLV9gr0FQH9SsowlrC6Ud0z
MHJLipXE+D62ly9dXnMo/zg+dSMt8shVK6IOd8nbZIQolqkEtLbGiIJOtcGyxF/SNIQV2UBPA/IT
290yT0DLExW9s+qsCPx9usSqXgMUZrsIA9B2+OCLHdX30sy5EJC78fZN+wRwRf5nmSS/YuW57Uxk
PQYavXQcj8g4u5EOf5SMKXF8H9+U+hiJRNMBskAhxaXH2HGFEiHmNrXACNi371F/sJsxiVYBcsDJ
x33QOUxGX1Ush6taZfYTA0dGpS8YD0G2pbaCvNQUCTP2rZTgXS8EmC0goLztrh6389CJ1zB95+eh
lQYxNBgt9FNJsgTk1B1f3r6O01vHpZLug0N0Nrytcdjk8mC0Fip5R3n838TtydJuWVNnbmS7H2dQ
QeiMsbELPstszMeTXETjztbRIgRf0CGd26d97UJRPJI5fDALtidlvszRI0TBeY/PfzrKEUiIYaBK
WC7nKKXdEpCut5aILv30Bgu3FwY8y0z2hXBTD28av/pJSN/ISj1AeAnZLa7doelWhFJWrtndRMku
LxOKmR/kQxWP3pndLVQFYgFy6rIi26YnvEiQimsxjtmEZU1+KXDuTTMMXiRIK1Oi+xNirPt44/Pi
5h2E0valshK1WFzZxa4+8JYIkCDhwvn2mZTPDnBStmfldzXNSLzMKPd0+//cmtUr1dvlpF+O46BS
yW6w8OPbOZIgcbRsbAmAYBtrl4AZbe+TnnESUWanPK5k90fK/rev/ETXHCk+Wv1sSeWAJ9qaceZe
l/U1ajWqkxQd+z8nwHGgoen4JfP+8AaWXex257b7lIWhRd2ac0USCt8YPm61Mo4Skua2DySVWNpx
gYQK1IUIldufhkuY90CrRJcUn/5yK1No+K2Z8YEFBebaT3xBOEUAk4t3QSk923zGpUnteyPyi2gm
fCmr6HENjUJFkT30ukOiMC7UC3X4TLctts2sFJAs2VvN/XUYpEzjST0R3rnw9+/sYJDJ+60lT35Z
HwQkgEm8iVlZQyLs2GjMyYjEzEuEuicnFyUEVqPAVPIhZjHvSh8d9IPavfTg1WDICElX1Cwt/6fS
2Ge8K/k3zwDsn4saztIiMlcpwScTo5zjKa1sEtPSOzJWgMrQOiAxRdWuhMUWuUI6L568emwAr4L/
xJQ4986AhKnUeW6w0RetCxvBf3JfNU26jvUE08NbDF3Jc66Ezr1HYsLJBxyiPB7BVLmu8L+j1G/Z
EkQf++Cfau/n1A+kJlM7Gj4XNXa4LA12mRF7k+0TfgVNQRrCrGLIblGo8mbuiZfnrlD2AiOSKvA3
WhIii736JOvgJ5iP9RssBa0uUG7LpJrtpNqhsW0gRu5gQEnFDX4/oX4ni2GiLafrSlR88mdpQ9wJ
ylw+FylfwSF1/joiEmzw3JK+Q22XLXfM3MRsA1TPjOq7FzzKbw8P+QkYPOkIPGdxq3kr8pBJoBry
s5dpYkjTATh/zcVHMHn8cl5FGQo3Du1oaUP9NLM8sRpD0vgymPhlXmfZQgpPvqTNuL/9ZNBQX+OJ
ylDxYJt9LKGZVhEznzf4/50A7tIzAHDRGioMp87qMLfnUL4O/3ToHo3pX8saznoNU1lf3vItX2ZD
6LnP5U6oxA89CJjAqBYQiQOvux3gYekG623T4CcN+B1ChWDlKSpdSCaExnQBDxRsjidi8qsbigF9
0KbPkHU/EfUdy+5wUle4IcvJQQTOdfmhqZVMpcEuxoa439085xHcQysiLQvWiQ5MJdVCQkUiscrC
4Wc0HmqzgBRnQCigSxjT363in4mib1ACU4h0fyOrSuD1eotRBqjZB8b06cy5oHx2lfFvadNJjyxW
GNsfK4V1H6pEWxsyUhOo966sFCIzhInNq8FpuxoFTKOJqrClUkOpD3u3JCJs5yVk9Bl9EsI/BIo5
dtXoVRjDHkyMvL0rPdCXgnjbMJbWW3QavAMZgPd2FNFnW6fkr3c6dcDUu+5anPoUme613ZTMWoof
nvvDIF/h1OI3ixIyqCej9oFdxphWkaJjnrn3uwLxBoz9DyWmY5z2rqOUn0pznoUrISkjfKkUevBC
j8BTZ/ExoteAWLOxEo3CMQBxVpLcSJZGda+Jn49ROAsLKGQtGizu6lo7y2NY5q1M4K4beD6W2/ve
PYsyYR3cv+S9dyueYSlmeAz4o+TdKDa5WvMLvHVCxBiM+ZOp7fDqVjiNSQmxmc0RLcgAPrPcfhXU
D0cJEzBb3ZbbQkXMxgovLXHL2Ud+HDryakEKrLsTYf232coqLiLgFyuIdkXOby86vqWhMknswi50
jz056ntxlVQ8J/hEmXZMZO392vuokJXlHJAad/q25iM8MKNxUmZFfEziV4Vx5c0uAm5si5qJTH3o
JlZHDjWFYjePfmmTv3gCInwhXbBkGI3GXqbmU4LwdRTOvSoxLV3vpqpcJnIqe2Q5XzoNvuh1mk77
BQCXVeguV+tsQTEo5g7Q5pp6/rs34MlmVfj3wjBZEyEn3MnYtZ2ddMRPltRAHdg8xF3DNQDuK1QF
KoFSnmtV5XkWBfjsPo7UXWDA05Ei6EQ7zA16vzv8YT47WaQg8ZwcSXnYa1K9T3mpCWq721CE3ck4
tx81zLFXZXaHN3w9jhpGszUzQfI1lU+80X5IfgpZ3CCSyQ+tYBwr1l+MmVindnqxjgodrvGjq7XT
ughglIpWAXoE1K8Ua1QI89ctJQaQTZC3s1EFBTopgNX4Lh9Z6FPHd/ic4JdxSGJJy/1jZa8zsIw9
eXkFPknRUlihVdQuKkau9w4mxAyKzptwekgriIASlenjKgpIBE9U/SazsStJrF4utSqkXaiJKfI3
WjRStVBY+qPcav8c+nK1M7fckmWM/pwsg76kL4UhzIOlBAEKuBCOB8C3fc/04+5eqoVO8Xq1P86L
rmBVgzNNb9uypQ4VqCjo+oGONhdo2U7n4fYdr7YumwNCMa1Kc/6f1Lz/4xAX7vo/2gGDlAYlKv5d
87Dsh6b5CnLc6Y1MCOhUmzgrBfei8sQDfI8PXriEJhrO89PVqk1CNI47UgCV5Wq9pow4adS9aWpg
QGrEdydaXThECkccOHFKJsaOJ97I3Zm8Ybt7AuO9SARR+4f+l0ZR556bxPN1rAcJd8S+fI4o3gkp
0y5+NdTbgh2tk7/X2M9KaXn/4XIIB0ZC6C96m+LfLrBAxd+CvvvyL6f39t60kb8ZDjC6CfyPlsJJ
oRhNRIoPA9GXCNOuBw2M2YM9vGNaQ0cBp5QUkUJdRfSOjGZ/2xlI6YjP3vGCPlzH2XLd3dYf8I3g
oBh16uOhUQKeCYZAEiP7+kAtWfDdIZOCJ9BBT4HxHgQP/kMbZ9MBGAiMbD9+9LmrrK+Jyg2a/ViU
0kx4jtjU3u03e7i8BYN6bQ9cbh7yhuoyhcWiptVOU+Bv0IDTKa493brSkAgD5bHv7IL9hpvhJDoy
7YnJhDqTxAfjVI2e4iL39lECFxd1ioJKe0hk/vtHJ6DovG+DfV7epcW4ITyBwHbIHCY9775Ws3FI
q1gMtW3+vSlawN409MZCYXMhRuZcdrQlD3ixuTzABAJjcoKJ/WgdS8rFcl3FpVJ8bw1k/A29t91o
LxE54LHZ+BrAxcTkkilABc+B7oqPlKkR6sjbsEVGO/XaY2SdT9RhMPTZZS2OvALfbth7JhdaT22x
tpdx77noEF277AKPEh4hUDeQsRHw/8GyZF53daNJBu5njw+ous+3FurePZmzogQoWQblB7Ru9ZYb
ya2RKZpYTa+Im1iSH/PncXbo8ugzO+yDaZvIYDBgG5Rf0C81auy5rE/acwQt8MbAiw3M9pUEJxEz
Bm55v37sAT7+slwr25TTKEqMvqnK6dvVu2mJqhRiiT0fvfcOW0/Is5BcFM8lc5vrDMyHzcWYSjv7
uK6Q2+6nQSb7D2VMyf/8D0Xbh0KAjPxFNKgE/twfLEfL96S9d0PImgtd5hUdA2njaCQv2oRRQBJB
0j29nC/zM9wL2MSFpRfs04HMCpYb86nnORNAPQvfubkD7NOj1lb8xCGnQnKqAeBSrMiWxREK/v/i
WZi8sAEcxaog623Xjxt+sxQLusItTFoHqXZ0C/mjbeOnntRP9pTrbeeGo8kkCqPFPl9D0gakYntW
Wy/wV28+xp3mQPgqOFAvHv4zyQubANIHWT40mGHPtJ2wcEF0XZ0bgtBSTZLoEro0dhzYISzND6TE
P7WdO6oZc0rkDUzGyAPE8BXGOVFNMk9cL7ZOCQhtO8C98Ya+PzNWmquQIwXXdK6e/j5MZMIPq9k4
ttNhzc8/ANvePgM9R7IKjDHbF990n1UgtolIo/bMMAYxz3+jOZibSCazw2xT4LV+337loBImPU2N
aqn0ugbgE1kRBtQfAHRr/oKcSjcQmo7k+O+8e+w4Q2TI+yfoZNtwNkPuKt5qlu7tuW8FNHdAgEYJ
VsdcwRiMcFAftwdCskGcxYQ7zY+iylflyQpMeD+8OcEnpPaxwHX1jZpi7AFxDR1bBJeHV/O+H9aL
/r/U/U7pWPKUghwFN5QTgCWJi7zDC/6zgZD29fvZdskaxga+OD5m1RvpZsySs9hW+Y8yO4nWhdLI
eOmFbf5NYm4ivWXqujxShcffplU+yJAeBWrJoGJUSG6Gp5+M8Y8OEavNX7V9r8T7JP6k+LDLVUVs
zZ0j9hOPg1m5cNlN9YgmRa1xXppO6/2SlTgPuNsQiw5ApgxQU/Js89dwpYqxa0Z5UX3CoB1UjSdf
l9JRwBt9PpTWj9yOSVx49f1J6cG1iexVami7IZqxe8CDbWW2F92I5in8TUpSYcsUkAsUFNCuDXik
5BSRw0EVR3APR13V6cJvhsQR6P0N5PiJeFnQJ+E3Be2p9Mc/2tkr1gerxAsJ29VoY3DdNDOA88qr
6z5kdV/gnshsTHFp9ubqd8QwKeau0wTS2MxeqW1JrkwTg+4GP0obfhbcjzmgxKIJGZ0Iu5Ougt9d
woa/32bW0GqJNky2PsokoQfP/IIkun62lR1O3xRu7r42U6Vyu7Z/9rMU7PbFTjCjBXgePPaa0bL7
7Q9vwL77PhoGV9uiE9MWZPOjpsqkaTtI4C2jid5NmVKvvhihQt6BFT1g+QAvIf/I5dWXZ9YE5HfH
a7l78XD8XiRDtYdKfvdimMD/STYkGWuV0E3C8GUdHIViguvXbVyVH/l01AwWyGiXdejKNiT3ae4J
VKTLJJsVPims+Cuy6V1kmyD5c5JxxiyL3MykS4P5ogWt5AzAj6N7WznV0ZVwEILOERAQ7SI4laLH
NsBEOTocygpAlbd/usxyztjfeS4W1mlO2f0r9b9nUIYkhhtcya2M6SyNEhYE9ERm1ppoBqhTsi/A
VD3AG8klSExRtMTw0PhLLLN7ngfMJac4vp+Uu0zwdad4Lq2VMCwrK7zPOkdEEmwP1J9pSqE7w7Q8
0ELdtWd6OfTJGyC6UjQiQtIqMWghjKoN2pVmNbDcYM14ghd2GrExNc+zs5atOGCnfMqGM9U2hi+a
vLPMAb6sLy/avGLnpcSfjlkDm5QjdlWIC9hYcqEbTO7t5TA+cr0yD6xFEgOTm95OsOe5nnYReg7C
N8KKvP5wIBdsgU8pOpayEJ/jybW1Q6GyvxSOX9S3bw4MV1mKEADhNrKqyX57zKJTRoW9GmyA9P1w
SDQ/An7ZxxzgZ16atCmoddwi0aUjCwg9YUSDWiyNxmC3CwEwKiEL6vtiy0nK7qeX+kVBIUZFdJcF
seIPYEFZzqaCa0kf15D1IHGfaqIXeHFK4xbbta3BWJGQ2UzXJ0eh7kNGosdWr1z0RG9mcubTzLyG
seGYemth84agAtiWhtVtI+i22gwwGOm9Wrxu+YdERsCYL1fF7fFanz+wIU+w9eShvp2c4eQdsAcv
XPJNdI0SPHatBmyi9yyI4kr5PdF6ZGtIMBW9kuxmPuy4I2ccJhIZpvAxiNXKx4uvh/21IRU3Ghap
sYM8b2kuzRCCFl5rHVY9DGr5UlRc+oB03hbQ3Sy5W8H11YaBqulP4MVmqsNGY+w9WjbjxJ/WZj6W
abdKE45e6jGuvaMcOb25BogRNT3ZszBTTlzPUKmzoCNc6drXGxtb2R0QKvR/IDrJ1mlPNDoavcLZ
Qc0EV8WfBN7ZmuJbNqHwxwIWGZNXj3YHyoLbIvTV4QmAYWqgQBxR/M0YTxzTqgr3DWVz/D+yApG/
KLbDqx/6WibeYhNOEoV6VwJ1eQEyHcMS36JfCcxyzlBpjTmFIxYTZsoAGUQ0ndPvGRKib4rhNrKb
0NMgZTRkpyA3J+Cq0oR+xFhpgxngbt3goh2kPYaAmQgbJE6z2PiOiir+EnAx8cM6aiJd8fZm9Q/s
vS+TOSivY8ofCNYW/1xekYVb0dgYtsjkk1aTaEf6pV1EzQnT9W4utX+kNtxPP4PuOexkUVeOUKXU
S3ZmTvYctlyfBn7sYLdlwophNjihBpn2hxMrs8ZtiE7oOw+wkXKpUSQwX7cj9VhK4gljdKkIuO6L
8sKvhg4MB+aqfQxvc/trZXmSpTKWGT/5NePH6emh9hBKkjYmKDt1d0sJshYjx20dRf++9W2iapy/
rw0iiO34hI5GZuyFSQlqAHTKDHjiuZjfC2kVUhKKFVcNihoYNBb5cU6Lx3wmhausr3mSIw8pWqu1
VNT6rpFybF463N9wkSQEQiCX641ZfHfdaozJcaCrREi2y3Ze9mkX53FUAKxF85JQLEnlOsEN8hEw
0xGBAik4Ed5ppSjKrQAP7ksovfEdGPKYs2YLRQAZJgscXMjh2qdi0xdyECw1VKp6yyZAZn9OTOXO
s0dx8aUX/QwAIQD71e9115YIzFM7xZtVlFi+Cv0aU6cgpkVT34i433c6PlVWs/wiZHKgNswRyS8v
TSLc+hYHxU3J4y0tWHrPEPI32NNXf4ndDRq2nvCqc6Lde9OwasgI4fpE85dpIeGQ769dujkdirMv
a+nEWfFvuhySkqmlB3ROjNF7/VU9QIjGE8IKNpb113orYxew8fOWyI2xVkhuSvM2V0418xCyjWkt
HN2ENZg35IBBaa4U2qkOmYlF+RjSMD0cLYEhYY0yHtvozhpD1m7CzrF7dQocmsXbP9fW8eHK+Ptv
eKVzKCVGlJXWp74MRaKIoICc6J9kRdEa823dhjF6PPmdDrRfpGgqYnbOH5xAb0l85NCf0OrZ5Een
LA5DiayWPzW9rmHEam+0uE1fki/GHqf5goQUXeQ6x/q2Q9TuOwGJElIjA6wUVJBuJ9X3IPGUgRsz
d6IOwRlEAsGsU9OJKmiJfkRfqmItcDZ/PqBWBfVKV1SAZBi131VYOVtcexf3Gv93k2Zt3ztgek26
tgQu+yxl6bnkMmIrNUymT6gVMOffjNKfIIiHgYFv21pJ5FHbPMROTxr1vBo2L2qbNXwhkCPYaF6G
4NFBGnHJoNwLYwnOcPMEPncD7XDVRcz9mSmvzPx0cPys7WdMFYCdr6UlBhZj63CUzNSEKXgNnDbX
cJOP2BZ6yObg0dU/kBMhwEL/J+lvELkKFqscmsbRcXK49W/J8DQ7TKlti5/Dqk9vUc0CnqPh54hJ
Q2II5tq8yA1AygZ3eowqs6kveO/X2r6SpzYIppzs8kchRm9e41GbI/70fxjwQEGnaNRUBCYolBE5
9SgeSlumfIkptJCzQiA8d2r1gxXb3gVj41G7rQbf5tOubucvWxsZiu1tB9101Xky7JNGIRSU3rj/
NNwHd1lAR+BpfJqSx3dQCWFJxqz1MG2RdSd7RXLNcSMjyMITOmNAys9iD0MDnmzJ35qzkmBRQSnr
ysgTibdRgGAIxDNhJEUk5QN7Q16e2aZo/YOFs7C31zVcYerTJZCDMPox4r3X9el7Cpgi5u8BpdFP
W4+l9eEVnoUPLVQB6kPCfco2oIcfuUecDvVIlTPFW70fYbI5NL714tENKF2kDRA3DXdmYhGyP2sA
w8bjteJ8A/pL+lWx4OiAulMcx2FmhoPWBs9qWwDB8V/BG0JDGWesj2LC3l0kVZd1d4xlLtZn3m2C
L43yqa7VljMyJ2Jkw5VOU4L2TlqNcl8fxh1WiqxknLl1Cmwjaco0KBbTL5MHFu1X73APquVXgkI8
Nr5tX8K8Cgb1vrHARRZ9fttKQKgwzXZ/prU4stepDRvOiEjkM+01b/PG7bZ3kIgGpbRMOxwHLf64
5MtNxMK8sTMBwpEM718GmO7wpMF9R1TQBxwDQjxIucOp0Ce4N3tC5qaSVG3JrRRDtWX7rxeqC2rg
7YDBDBdU1WKyrI4GppCyV5uKfvLDYnFjuiCBk0kmecZOUt2blQ/S2UHDcBCf9myLn0oFzhCrhhHu
Xq2+vjqrF6BbsCRlq90smqaeJFWzfDLFoDqaRgNF2TChT4CNCUyALd9YEuUyBhSfMPECyBnbiUHm
OMW7V1qELX4ieJs2pv77LMjmEQEMsX5/1NVocivvnbQrukEtManB1iw7H3Cap7q1YxJSwBLz2WHR
CbTAx/9yBchELnPHsGz4lulufhkkUVSItVwiRYKesjLqQA0IC6A3Z6Eaw0DobzOWH5Eg0e8bM527
asV5XokdJQ8eiGzqT4dbIaxXqSJ7JDvx4JeGc/AomK8nqDXMF0fLNZYws9XBHCGuZQR4nTLjsujH
OZg8BR3DviSFOhX3F7HZAZJYda1CSlHVU3j1hCStPb/b6ezcVAGA1t/t6AXYkKm/+eoFwyoiIryf
8zYk8jpKJZfnopxgQSzoYlJsytv4Q6pz4K8Wuhmj4YuFyOmuMURriQom+DD63drf6nAZUTbF2pbD
oiUlY9wdE4SRHjhdHOn0Sbg4IzNfN/Ufv7zeApFOC+fzJWK2Rd8lnBQJ5qh47tTVBGDbsoYrJhd6
GnXQ0UkVDkOnAT8MGBZ+w4W6dUZZT+3idZonXdgF1wKDehRtMNYUz4VFjZtViDFl+XGZBW6HLWJd
M4ivpV7jMbN0bRjGlKm/Q3kwS+QCk8ddrBULUMdU6reW8ITrCNgbw0b/Kl8/sprbUV5STNVZqrSE
fAl9iWTtleGVDAzFTooL34+n5mwcFWf/b1j6f+06mEOlbtH2ndOoeUbOt7+DLJbtQWnCxtxKO28Q
Oj0S0KLcLtLHpNDXgbKBaoyW+LaYol+yCUbb8bWvl68UqJIX04beGfbGtXqIBE8PzmEQNl8yAlqJ
Dx8+0555IvNirYQ5kZ2rd2ehIo7pQjA9d1SMGe8i7j2+F+zw7VxhPQjfZOcb/iQWRQ1pCZWOf3Sj
VnOxqDuvD6g1YMytC8GcI9VYi1hKyoACoduWT2tsJ1kcX6yCrJQSOMArS1EOvsR0x2j9QXQnURxm
mutD/ammImGLLzZKwKse7G0CMHLdZUFlFmZ31uscR5jB+u4B3Hd9LxThVuaGMpV5TgG8UbNziFBA
OezPDcz3l93e/1A6oXezRK1ulog3bus1ge72Ds9prZxzSibtq3mhmTJnET9loEyxEbkgP1SUFyBZ
eBBVlQpnSArnaKxZL/1s5Gl/l6WNix01sOaWvBQyAxd3GDk/jQf4fC+bK9dl8i+adz81atp7XNGX
f8WcmKA2+tRw35jYu9zBv0KaaLxoMlvShTlOxTPU9zi/HZwF4jRwb1g5z8r+IffIOgG/4QN7L49c
tO3w3yV4Deb/xCdhaP+eha9t2nhFmAes2IRyG/j1O+xiDHOquHoAH7hH/QKnC7A8di1XOMIsRFgU
tsXC3ZGZFPbCFio0GpsoHJjxwLqDk2h1GoxjPFR34q18AZBH/zotpv6T9yiVXs8xLyPCGP0gtsdJ
djPPDKYI49R+JkSmFMHfJx2KL2MxW4ncMbrL67sUYbpTE74DNwhcimj12bwrPdT8RMCb5omdEUxK
MHTSDHGQp62xUjz9+KRJz91w2fpXSMOlQgaSglaF1tVaAV8aZRFIY+2Ngnq2ia9u6PSiYogm+1Uj
sFKFJDwkER5+r8Hth3oV9TriUPE3gbdXwr9+u3AbsqrKzQCYIHGaS7QXaj2GdYv6JXyyCwR3IgCj
ycUQHjA3rTGn/8rNi6fGynw3pIHQAlxnpQsGVGYpuSOmfq5bTOiFt/VxzYqC8bxSttAqX7VqNLc+
MloFCQBUIdKmOAo/2EAIFr9ADnAGZ43DwhQKS/egzQVVJtjV0Er4zOmo26v6thcanu0azAtcdtKo
RWzELfeITT+34p4iWKy+vAAHEYcrDnZwwnX2+aSGOXVhWu8+fU0Sw7EwHW5K18lObTxdxkWdCfSt
jhZY9uvGHyYIPIULJKinxG2Ttympcs7Bwnx45Af+FBwsPQnm93f3aLRgFgqRcBjsVw4gG1KyGvna
nXG4KtERO2oXcVeQPZzSYrWY264EPmAk8ay/ye4/6OZ7XT8S1gYuF1YU/cL8Oon5nWZ51qCiIm1W
NyKl0GFI43EeKZXw5INA2ZiLBEGyLkFks8EeC2TJCYUEwc5JFA97t6esEGXgi21PtM3I0rS/jU0k
MTse11dZbI81pQ/tUmiXO0HNT2GGFVNeO0rURAlmb0LWp84ufuAppKGXdLZECV+tO/9Ctl/JLzMD
pDyhU5bjyD/1NoFT17OcQahFreqcVMutATHWSrldOQEaGqsLMS9Cwd8T6eM8zTXAJ02JGcSx07Cn
AKPyZqPzkKOIIraHUwNsl6SfvBnzxOktce+j7EPDOstjfU8aiKiqAFEdvOah0S0qpzXoMSv0y7JZ
VRBszoxS0XiAxvt7FbgMxFcIKxpxW5nKaTFfxhRA/ERQPg656kr72vjV4h/bPeQycYdRpAknvnhG
4S5VDIZCxgNn68F7NYOraR/e2vvLyi1jlw7/kkddwT+IJkzHJRtnzKER3Ovq3n/HY3bXJN+8fnDw
+4Qyckm1kXVQkqLsFM1ithewf4iWlYDg9rQ18JF9k1+uzKxlM3lIwYrcKBLDVvEYzoPi0GvHr6Ca
WcygpaQIHzDufamMBWmp932iOdCfgtXL88/fx+RW+4kk7tTYMr0CQjpRw5JBIhzaS20bwwQohsvc
awUfKdVjtnOSoQLn6n+qx7gRHi+CR9ULTBhs1tFPNPRPKHG/yJiy5m/YZZWatUIIhHca4DD4B7xQ
IO0s61BHkfFPtCEKJpPSxhGIQd/x5+3+679dQCYQ4VB1ICNJkYHO96zMr+nIXhBQMNi+uUoQjGJF
10YdsXhpzTFGpVrI7bZN+y/wAglJjM3G4GJ9v9NbUPML3TQMNpjgRKFSOKpNdtcBA2gy1Z5IF8IP
avx+gujoHZz8+j9VDgUIk/8iYn6tofEEmKPVquAiOYhOlaJO7mymdw0mpgQ4n4zX+xE1o/Zrnxse
fzinhPcFgGHvVQPGvjEfxFki9RC+xEW//QFtJ9T8u55/3moZ+Spsg0FrBCDvI0iseLQYK4/MIkhj
aoCfyawX9i68VfKqT9vh3StxgvJara++ORMIGVlf3MpecPZZpagwnnAXVUJeC+kKPkm5IHCWFM84
jptjaFV+1iZnmzeTGUv5V+F7GMDdoFr/e53HSoifKEsocmNwowH79VL5ypTTfjCXUrb//ZhtHF45
z+zAQSxMXJFJCKBe/aygV99JByVLnPADl5glvZkxb8G16d6uDJlS1UsIIDITdJzxScdMiHSYr792
S0iE3mgL9buDZCS0g9WhV4Bw3EOLzfIorEe5adTubdQWCk2S1CDoaLV9voW25pW8sLe3yzrbKElb
YmLYESuS4Q1UvvKsrVzZhM3X92wBG6c6U9iHpVnIJIElG9960vYF3RPuCwIDMsfpDpnDmKU0KsdQ
JJcFpg++6ETbkLsHQhgjT2HlyqherQp4hnzU3EQX4SGf7I2t0LBvpqCNP0fffglgXxLhmx3ADnWy
qyJPsHesF46Pjg4JF96qL3H1vt5ydJV2WfkwOMiZw0lerNjR1XRgggE8eBzTmor9YiYWT/DUHqx7
aKwOoAXP+us4JML0+hEgIpAE2xenMInADOih1ka4vQ5uHOeMIdgLUPBSJgVH2Lc95O19mxbCES+K
b+JKqgwLGs8Btc4ivi8d5/KHW771rCU/jmIrplindIKDRTOuRhz5HKSer4F1+eSelvD885OlFqZN
fzloGlPvLE3UaHkhw/arCyVSdYVs5TZ54olWFOgtgZpzKn6ygsctwvv1h7K/bSSribTmQXAhaFSd
Bbgg6brVVa0qfiS/TQeFCkhrSgOK/w4TuRuEekLjJYC6zyicCFAmRs0f4voHwkDl0Dqqlaj6SRDS
57h2yPwCIoYsAMp/iULZ8UO0mdIwTbez1isjmwe6y4PgEfUk9Xdt19H7nOWAM0kkj/SkzD8ssCWb
naMqP71kZQAnhL3Ivho5PedIaEYjKgd0GPgDUjH7eHwsX5onKInJjRZioO/9qwkEittwml0y+8Id
Zi61K4/PvyKBhKAHnzWQCdLL85Fe1BN6x38TPs7lZVjw5kBna3cCoGrVpEGyiZrcmPorT1aP6V9E
UfWi6hun+ZMFjyVTGS9KsanKo0ZhS1EcYNeqNkxSeYse6emQL9HCyRqZayuvIOyZdGO9+kJ0lz30
9PFhScic0JXpoZYH+64haBp41GTzl+fZ4Xoh3ehjPKO3NpFls4IIxTOIqQUBRvR4JjeP439hEfjU
MzHv/NWlTlwF2bcdkWDBwMe/0Gq2DcSzVA9mLiNYkFwlq1T2HmNwaW4XsCDS3I0uMl0aAkUXl8Xk
SFNrl/uwDvZFfRyk7W95a4kebKvoZGY3LyQqJjZ/eTf1NRhulEXox3TeA1aqqhge1hjJiDf03zvL
am9/A5NLJNpcoE11i1nzzI59sK8RMN2xsxwoXBoW62kc/S4m5OsGRu8n7jVZPvV+/ae38hM6lQcV
xTFI4ii8cDXbUaQEcZ5zMmF6RyREh6KXumN0+zHng2pn4ROHsYLaNJn+b6ocLykfUGDJCUJx6FaW
NknTNr1MSF9S5v6JqMfT3lb5hc/jaz0j2df2Q1VlhMFdBZ4y3Z6XqTsurPvcchp7PBqY/6rWImLO
DRBpTeYNLEm7TNzmgyVyBqD5OFhd6FnmINNgsrg24XsCJO/uYNIo3a7OYxj7WCDN901qsYu9lf8b
Ih5Wb8l6N8P09pA8sRBslHXu0ULOK/GW3P6C7/mlVIjuINMeMHCOzAQcl5lv0a0pz4gNOVe/fNbO
ikGUKNbnvPAAOW8kBbsZVzv2hgz+HKHAAEGhXXFxfVMjphetOk2sf2JhAY35YwTsiXLqRXKCjq/V
o4C0XM+TYt+SwCXdJsz0FuHr/GVTLf4jmLqr6DcOHE7KZP3cQwr/8h0p+Yw2HpVBJ+cCiPqEyHj3
RmGIOkYq3DtXw8gvr9ZWYcSvHJZACVABAT0nxSnDyYx2nCxy7ADyIl5kzQjNZtrqNNaERE0OSihp
EHJU6EoDEI3qBRvhXtee4YmmQ31Zg3nH79aDcATmVWDqWhg+yM5KzmaQhZu6W9PU798AE5VpG+7c
o3G4A8csw+bFy5Om2K/OJUgoVae1Sc0KIKYa7T+2DuGqmiR2v6q25I66/AuwyD+VE9rWrZ8iuNdF
K6+LXvZynJd40ED1Hc5S1NG2QhC++OC5ns52NmM47ZqseV+Jr1pgnltkZZ6LaZe14ypRh5xf15F9
kGoL3RpB+1P6AFNIPtgSi3UzkPDM8bts0YiveahXi3V5CQdqGKbD5yhmd5sTO9UdyhCIXismnMf9
ItVTphCuuGRAuEbvDeZ2vfXrp238vkkVZ5B8t369l438LOf4/FuLibixU4zlHpM9AnVxABu9eYYY
gziZhqw8xlU9+JT6SvKsV2UO2ElaUPgfogSPWPTjoHauOlKnKPPG2jjeFmTzhSZGwYOM1YU5jAzn
Ba0T02RaWSiKgXxdfMQbtZ50O6pqVLCUUs6mUt9/aUxTcx0M5FPbn114nKrSFJg/UIthKl7P2fJY
Gii8MrQMiHNRpylmazNQl5OoR33fKjCtC9UvaGgGmlBwik8DBFrlKduVgcl8AE2nj4kt/FHGAPQu
FZKYliwknew/ZePwcZk+Sf5zZH8f+8XOBeTJSWrl+Sz0Av3LdXPfWfi0s/+df4YVtR4A4eSR+lPI
JCcrRe32SQ6RBmR0MbGQS4y/vrQG6b5JNBOsx1ZWPpIgOp9fTFX+G9WTNQRW6ngF1ZLpmTrcDUUo
A928qfnKTeGE97FNjlz3ANNXNXWDD5edIKKNi3MezjwAuflrKYu3b71QrlDN9fV9Zhrwd9oFNTRL
VtYca9uR3YzaJsHgS0X0mo504CnJ6DWxd+10wnmN4Q41xMQJdTjLNHqvbfjRNjBdxz6s5lalpw4u
nNEHXBmu9GyV4lEuPbrj2Pc7n+10f2cqNeuIAtgstraS8fVDxkwhcS0Tca8/QX9wA8Z/CxuDUOor
khfo8FpRDZu+7jzMB6y7A6dN5HXQwSOfKNyvdM+tcbSIyLqQFD++FBA/ryzzjw0nhBEYz1PnLAft
xY4NJAFFjRqWw2TNrStUNUEzbo/OZ0dPTeUDxzxrp3YimqYljGBqmusQBu3rn8WrYXGzak/3OcOp
tSEArf4oARqComQ3v4nKyr2my8PvnAUDfW03ioHxJsVWbTptOMPQiCO9cxgYIldvvA3ma3eRBBeR
3bxBJtQDgQSm/r1f9nhrs/QaZo9s74XJnlzgMBnUUbp77R8PlAppGTWh+REqcmtEQ0oy8eLSMl+U
ONtdzkLRGm4CZKBXGxORBxTQBZBRMzYyDOjWwIxaTmiTTbulVeqBj54vemUfFQ18fU9kqXwp64uA
7Ozry6sz5QWWzgg0TbLMAMwihlOqJ9knPYlUiNhyVGKgK0q0KeXhbBZoyP+NzGN7RPoQhdSJtHMv
43xUl1fuW+ZBLb0ELTl180TvMc4WkujI3/Yz/eALebAgQ1/JGZBk3kskriWTKnaPrfS/TBXKvrrw
fpR+cMRr56nj25w6viy1bQFX3oE5XVZ6vPQQXQFMf2aQs18K1dMn3d8MTsi9zqVvxgTBVJ5vNapu
ZWap+S2tkcyYMhFFOiFbNqCXR3WJQpyIdahg4rgIbhlEvQuvg9phJDXGFgPGS0qAtptcsXk0XeeQ
/RJZng2BqJ4aeKGKpXhXIclNpm36Ir2j3TMjREKmXQ/SrKs3W2MDMueF+icTXSnROI0yG/mnEqZ5
C3lNAmS7SOKiiN9WEQUDXJ6TL4ttVR08iu51CxZgdnVtVfkkb87FHDZh4PTB+mLbMNMg6ASGFuJO
Zi8Swa6EHKLoQpsXrYzXDClXELaVk9PLH4fUbaw4d7p961TMbRIdknmuVWcgEJNGfhZQ64jqoNEL
MKdMdQGhFRRR0XrpU5lFtD7ne0LwmabjTbtU24Ic0DBViw2UASGwGJM4dxu6gjOF6IUI/e2FgVdG
6xLCXu0/ooq01I06MZUzy4e/YgAF7pV9JXnIozPWlWYUPuWZXkrIOnBw85hYxRZeRRz/G0COT/6j
9YLu1HQMqzkmwi22Bh7UjUvzC/r3anasZOLDGN5ZTlTGC8sl/KWHYaeyueSvAG7Ov0yXZi38aZdg
xn76P2vmql99bA7uDeHIiRHtj4+dgtQQ0WK+u7UgoDzh4n7k+2GvKTGtwwdZQdeKaGpeKkwrfftB
1JduY70i56zKFsUF7LB6WNfF3oejJPl8bzsBfO+hF5u3TJU11F3HqLCSeyPhOtfPZEsnJ1r3PSUk
BGm7s5zvM/tQvJdIFdUwtnTIQV/z+XWatGKwe7a9M5XQAcesXclQeA0M1cma3hJIds3/+hltKIra
1Y9aHpYVdTwjA0Q/IlzHBBxFmmF8YnrHXQZlT56LAhSr/7ySYlrnkF7743gLi4O6ztG61BKqQHbV
gSu3SrLzR4PMuXrNUVjTB5/El0cqAcMVEwFjBxNhq1tmOP8f5M4BfurSaCIP1KskCqsWM/gDv05Z
R8o09wkWQ/IP1aX4Hq82xnt0Ef6NiqQRCH+z4k4QzBdKbhIZz7w28dY0FLPdDRonwAJ9M9uNwg8g
fQ+ghC/tMQTD/nxe5ahdz+6PdQkeexwd0oQqKq+qyn6XX03YSVJM7UixLpOY3Ul+Cd9+RJ8sdjYc
bp3Cai3QZZ/aFuCxm58z2TBZOOibZFdQgZAhISt3LGgr7sDdsw/M7xb66hPUwhGtk5PkYlLa1ACv
7dETdl2nybzqwuTYq3e7+GZN4MNxW6dfkgXHGyXwfLOYAAgNeTEQTnfsJnFbMJ2+kkeuY6o7jdvV
MWJR27qDv27KTI1TnBoG76/Hfr1SDBCIn05CkWAa+dvC3ANyn7pV94F0MNNczSZmQus3uQsq7pgh
ZGYJr3I4bfoxtt5vt/J3DoiAwFVVjmGK+LeI27IX9MF8bZRpJee9MjoRUVhk0E1LaOVXoIv6bDsU
L76rMK0Avf+U6lctBdTYkgo3IbTKMQ7t1tK4rRWaZ+i0pxdY1znIzkEc2t/pePIh3I6jCcjOzj8b
e27wUA1nMJonGjEIgH4PIxkNVVzADhrDW4QI2guDPSkSrP2j6LCQ2+reWsk3JI4if5gshIQeYrnM
/LdkkxqlHmNVFOWxcUNMYXSD6WCRcVanMsg1Se4QSUhNvpeeDNRIXmJf+JWfsu85xSttkd6dghd+
E9Y0utHiIr0rP0dAo1fWkHHgVs0DhHK3futlBzAkCWnKvOkwOTpbmwLo2smQynrxufswumR5G+lR
xMkWeN62nvuSfoZHAh/JYXnBUv2Oait11Gx2jKggz2qJdtEH/YOnU8Q5H/m2QWHdMJZDp2PXujtm
rAfyjkgXP0ZBSe1/wvZ6yg0EXlaP9Cci3KscyUAU+0hNtWR2Bjs3aqAnhDWh9NDnl0UMjLX4rjQS
swA/veAkvipUh8+ism8SSjGQ7DrsJ0OUr+qSEhtLWWfTIpTyq2hVUmz5vggf6NZITt4JOaQItuvj
BRfQuMt6H4jyW9XUC4uVcHIsMBGCPNVEIPB47F1vuIiYuGxie4+XYoFUbds0uFtk325LOEJ/Eire
NnpFXQbaxXIII2HwNBzIIPWWY2cz8CZCSYdTa4E3nVZP/L2XncUjeSEFjOZKFlB8tZFn2UwvRxUv
dJ4v8ZxN5KVMcmIIHiG6obHBYXQqwoZ8Ivz7suFsJjOXyAELq/rAF488Xj9229GcTHaom3ZATUWC
S57kviCw1WQMSx1Gw8OsPrOGDBq3AKCmDyLGtBB/LELP6E8EWVPqzOPv2lInv4tWctYVUeoL4fM+
yK5hmkht1eYDOgfPh1VUoNGgj4swXN5QyGr+0hxcTG3ny97czoLFYM3tCHwmUQA9AbL8l++A46/y
5N8i0NuOFe6ovhPdGHkTKjaPhQEW+0wNuaYRmNQqpGf+CB9GuH6cBmXygK9qiLfB7knUAAcsVeWL
vQukQUSL7hssGVJsjf8uoWo9m8rmyLwCYeotuNJXCKOyHYCpRSt6gL2k6Y+CHjWN5gcbAUgIgUHJ
7ATy0WH6VS39Ck5AWiOhrpjfnbFLPclLI0gQvHX2U8LXPq+JOArA8DydLXZhxap8pAq38g6hgsZH
gVZIVAmC6+itp+nPL5MX6f4auIdG85426arHWt3r8SU2K4ngEWqs8awLMq7kauEFCocA1UYs23eI
TPQHGLm9iYk+nGTvNpVSUIXgqy5WxJYcNzdhVHdS+ueo5lIjxyB+xkGkeRMStmOvqLp84P8A2dh5
yuBP50k3T/+y8TcXfWVLvPTX7BEwpgrk3YvZINhK6CKekkZyJgLvgx1OVFJNkAcheWKBJzDSpjW+
qigPkzDwX5i0b/lU71THIti5Px6bHtaAGOL/BIEbCv5pibBsqA/FsWnrQXCH9UWTYqlAg47CrnzM
YOGReQ0jEA+rf5IuFUG95CV9m5XHDGAF6Dh8qUGrFG7MNkCnqXWIRi6R+/9Q/eOy8+60FIHvkgj/
3KgeeWcvHgoFzFBSzQIjuboWXUy5q0OlBkixapSrCTtoneLUTo1IJUT9oR00KPVD4ngfnZpCWpOs
H00n/a920xw5D1jVug23sMPcitle5OvKCvfefjzfG30AUySNURKwptoqW22Pk/vuwhSW0mcTmg/O
BIFyPtP1LmrVeYB7F6YxYA203et1UDq55ZFNkSzWAajMmN3P3R394AI7QT1220rkvN7bRODFr9Yw
BKqVa+30LNinCkikRb30nlYNsCT2bq1N0/qEmEws1aJ28eGMk2UkfmFjEcFtu0lG4gxZUpXRimw5
HhBbYrXZrJEDkwSQIuOsrtBjFuWOs0mhIWPoNbFXlIjO5QcrNKB2x3Cq/C2RRFavBJFuMPIbAnGQ
0E4TmxTAqOoTXWDum8bm19WgPTeNjkMHQAqmEXqcia4b6f/xOLtzKWOH5T/ZuTM5mDq4fJE01F1e
P8Hu0aOTH6c3s8+Y+DKxOj3S+zlxF//0+xiWpfGoQrlCXpeHRQdlR9sGAcCETfcS6aGtqah21Zxj
Ev8xLL9iaPtEBi/uyeqNF189ZAv2/GQZzc19rC2p+Dp3tb4JVCIiqFpPSK9H+veIncPEnfJ9QmzG
h3YK5zZMdK/v27Arfx5+F3dRw7NFYi8EHMshSHB9cC4VXJxbM3N8WZW4sNzA16gH1QV8v09HlCeM
S3kAtg/dQ9zVtJ2dVcnomH3TdQB7jIi+Fl1ZGD3OGSMX9LZ1lSzK3wKGvJ2s380GN1smCOj7M5UH
JKtdyunwxF+5zjSTpJ9dm0YNxeh3fpIny8slojphD4qeInLzwzq5krr0AhgbacvrzDcoB6f8UPuq
6AOGKEzjxScVgwYF8Vpmr5f0FYsVArv8zOG3ETb3MExRQFmCQA/lt9f+NuRHLj8bZhZEKOZecOlA
BM9pOtrQe32UdtHqK5iP8646f9lbmXyvbli3n9wPzUbIxRdzrYRHlBA4M0UCa1C19fl22QJlEmzJ
yWP5bjMWYNRLZBF8lOtTvGPAqGWmUYBFlv38KWIxbeSONpWM7BP+QMBrE8bEhrj6XhjGwGBNvQyn
Kb5uSfWkX0424sD2UhTF+hexrH+L0alLeVEXT3FggUG1UFXVDiagz1ZNOPWHtGw1XMl8ymZjshhJ
PyzMZjLbRD10E8wADywYB7dik64OYPZtiLHXtWaRuCObw7hUKKAbv6JZlXvGtvi95a+b1RVvJKRD
8pF/byflL0gO6fBvLgBmg7Mq6dasJm+xjCzxiJPHJlW26QN4nCxep3uybWppjH7oduVnFF/WuhfU
4iZ1A9FTMNDKPYbnxul2nHseZlnnfkKLckz7fUtcwbnfkqKUB/9sZ/wrUJOAojyhmhidTWbEsfS1
7U0lGThG9eG+h8yPrKve8Ajda2mTgRy9Hiwfg0EOBV1d8v/8BuqE9Efb+nrBS4zBbHRweSzARQDZ
PswNvAnBYl/UVrl9tDanN7o1f4ZdRpkC2bBzTafIuTZWTVmBvqRbhh2RxxikI2ycABjsIcoPULe8
Lzx2DuNxtJoBXrcv7bpb51xbZ2NcYEUagn6026qntfJON5S9OmGOE7ck2riXp9DCqgmaExM0czkI
V13DjeSHdlJxQpp35Li5ROVmrciMaSdOpockFU897iP9cZT4VyU6DW8ZCkifTfvFNDFl8cqvFWti
l/AbSKjOAURtBxQoXaZeVkthjCTrsQHEjA7oPPF9WLl5ey7qz9w4hZKVdwPUMbdjAY65qiBBH+VY
gheqYive/NSJz4ggSAAoMYfP5XEez4s45EG2g26hXUFvfmv9xjoOLCxVezngbtakt35FpEd9+MkD
1woSnhvmnt3/RrnCVao8Pc9IIgawo8jd8X5QAAn3PCd6B8Sd9sLb00564+D5LAX6PY4x92scVKOB
eFAm0Pi77OOuG0mZBYU7IisYGaYwm1Xos1RzNwac7hkt9k+YR1/0TSN4jeqjca7SY3ExA89BCtfy
djq6U8iSS7vvMYqElaRVeMESQ108doiFQBgKWkadxJhBwTIoCPF7DPPI9O5DW3vHuOMtbksdOL7O
O/ZJS77JXNVNSwnRl5qB4Lin8KEtrmtheRNTQsCqcLRyTs1xslyiOV0+aup70eArIsInuacCp8Qa
XkGHe0vXcYpS6c3ZK8MtQRlDQneDdVFOTYTJ4UGDi+4IDTjAMovNeNLA1m71STSrH7H+TFoayqIA
R64daowbxv4PpjdX4uZditrmdrhppwEi4nGTYJcIfOSJptxnd/vlBoPIyffB8+WIj7db1Jjeoocz
zlLJ0X0pdEgjZ3SWK0iQMGPfmAI3CrFDnLjomKzCvIVYJuW4u/E4rl7vQAhxApHkZMUmRLKzVlj6
Obyufbbiy6/CW9oUIN5h0dCQyYM3hm18EdJI6QMU381fy/56/4F7cgrK/4vPtoI/DizgtgS8h92l
mASplkmqufqR6xW5ikxWTACnM6g5qvwzJL91PmRQfXACW5V0UC1ewWC0c7/VAv3w1tSBWjnmXcDq
+hLgeeqRrzFX4Jsdm21Mwwioh9YOeQuzdYHaqXfZzgHeRqGFrmAncKl74XhLiKDLApFKqi3lUH1T
bT2Ynx+xap57DyBOKn6k/TQa9lakKx6tDHor8MhUGBy9kfplciZQRsBw7Jl7qx8P2WU9Rm5WG2Es
TN1oTqOjVTedXwEGbQWFyfOH+JREENOw+zS9XBiJHfhO2bQT+sCPFVYV8YCsvlbY98AszXNUzuRC
v/3qo7/NEQ75qzBVkCx7Hn2hQxgt1f/JmRFdGWg7KKBK7euRDICVcScBKgzHfluSWaPM/eXDOTTg
jH+5WaBTboTgK+PkvDd9QYVvGAWBR4EhjT/du8sqwABJpahtFi/ZfP3QoTFoSzS7nqN27hewZxBi
C/bNmqKyQARzqjfPFSOc2IXwgnE/g9eoF4dLIlOxYR8OD6VeIOME/rUuGLjqlblOdc5AQNZgTr2N
qx5y3KmUd8WOyskabLTTLPflz5IgD2iZnKZh4fTjAHub3CHIP1ocjvbMAwpvQJT+SclVw0kKJPfV
0RM6mTg+I5RO1GwQv8OpaWHIAjfyrTn9ed+NU8EJpZh+4g1jfPEHH5C6EZixjfJgPKHyrwgj+oWs
EyMEjbqY112ls0YLGeEM2+5RT/h4dKL/2U/Nlq6GsSI8lX+LY8A9Gixul2IDLlX7vpoWQY2I+Azy
5S0L8Gk9rkp+T2kdfxDn736HMOU60gLX0bM9NdI3jIgNxs34FeFFWOADK+xMaBB0+Cp725e51uy9
j4LMcaweget7s9yDmIyE2R+Yt85FTDU89JiOMeeF06N7TzXeZryLdOElMwM5TxXpBwvy0CdpXDaZ
dVkMAyimJGB1J8w7pPfbPp0tZsKF5mFoUmDgojzuo9h9OSNeQOo3+s1lOIXwbIEzNP+oewCsd8Y9
KPALOuAxBI1bDdE8BffYoIrWXqMKoWtozi/Puh2BS9dqTI95cslnQaYpDD8BGQoElNkzUVuLAJIX
65pitcqYLfjRF/1p+ELZHDg4ezY5e2rK0TMw4M+W39hg34ajDr/4wx16F2W3uVR3LBiuIOep5fYp
3Xq2EdFUyo6KRF1C+GYeZoboNK1fVGE5t0fTbypSu1hzuajVP3pb0MoFoN+wbAvLw0B9irDDnoJL
+ZASfp8z8E9dwgzYG4gIdXtYWXNbx6blPEM94hyf58mDDJ2e+CoPyhZ+NVt2tndg3oGzonjmVRWJ
jLA+xIkdOB+O8Q6/qPIxVJU5L52fC+4nmP8HRui/XfERQDDorZOSFyQAKFCvzwh98ujez8bkNaIA
V+3tViQoT5bij9jQXAu9z/mRdNJvSEqvPWNHL79Fq0kCEuo7q6WiYdGIYKGBcZUao1BjhmVYQvxI
VzSr1BVT6tPFqdAFsnws0MM9y8pqY8KLzikQlinAqdyqImoG+lgex+NNaj0zcz1ZKAxEY3ZQNoVo
h0J6WuDpbwp3SBARQCpei+NADFeuIVE8Tw9z5Bk3yjFbV7yR4RfijTS8gZGBwgCjpQb/qF1jaHyE
0en+o933Cc5G1+rCMp7dKROs/dM43qs6TqLn9YzLCFVRR9TNwh/hGt1rPU5aDwiqzVFX2TEJWcuC
A/ZlEiONKAsRRez3BYPMIAoHHWso9ac3ijykeTRWqalDx9FPa+1VUpZTMXog0EUh5H2r62/MvC0z
HjouTCyIJ8dM0PTShwjUeCkqFYNnxtb9lN9Noe/So2vb3mXwnNaLmPTlK2sf6WtkIUbeBQm7kZGv
vPCBQx3qVWy5ZqfFpohfeLIO5/DBS2WZejXG1XDUxPl0adn8WFBVnCSKUs7Z4vR+k2aEjBgqudxG
yTo0pif1kz1CCBGGGHY3tnKxvIiLvLOMBvGY2XF6V8eZzX4v+6nFrkkiesPodW+G3gtA/lbXjRER
aL2BUATeVIdAeqVUu61mFeYXRD99gqL91C0MkT44+YCX7bI50/eNI7+2rTfzY6tlyakpKJ6MQzwx
ZK+lNbKCJdzGpyQWXkEpaWhafoiJxCtELGxXoCS4PjsRqUEjbeQu780mbDFIe6sMBC0bO0PoaXBP
16G+G8YZE37AKIR5RTIU3anah6kfc91qmbwio90Fi1FrEvfh+Lg2YoG2PzopXRmDc14pjihU+RmF
rJmc9gq3xcsMl1gEi+1ZOoG5fYECfDfMiivedeOMdvaxIGPBTqPW82YfBFmRbfAjLiDdZA3ZKBTr
IVrfamCWW4qr7FwZ/d+RI3pWmkawTHgNAdHc7qOgU0yJHySpG7uXKmLV+v/xBqLT52SNUAfM198y
qRDfbDfFJa7uIhJzAkv135jhWNEJ2l/Hwrz69xmI3N0Mo2foemohk5v9bDYnYI7K1Ry16/A5ylLC
no9Dg7MsCvGsDgCyTq6C29Wuk1RDB8a+MvHMsnfHlpJiTiDvM9KByyJRZA4OaC6xG8xyIxQL8X0B
jsXx7UZGUbgiqVIRVYC2XT04EVoXahcgn1qoh3FR0kMLtMiiyA2GGXipZ3jQ5Go609rUAX5vMwe4
K97go5PEPRk5UKuQ+bF1nFrs5mr1RQU+oM/jB+qERe117dYSGwLFf8c9r9Lag3+l0nA812b1Ve57
NGuIE5zwylIddrHRQSTab3NX02nhO0+3h9hs6sEm5/7W7Pi67hfdOsWSRBYRKQ+BjlTwesaHzvtX
dutu+QTOwqq9hvek3sH8shjT6VsHEvrEe4uA7NjmOpj/2OkEyjGgaEGv9tnSrF6sf89N4N6hvvZo
x9zQ1AnA4qecOoMw5ZJW/6rcTUob+O16rDhzNgpZOWG0m8KeXOXkrtXkJY+QpE3x4Yw5iRTV8nUJ
DnVWxEaaamE9PdEq2jKoX++8xgXpD/FmeeXdTHJLOcfJGtrsiFFC/7teWH9CAJiF2FwmF8ofemEr
Of/S7wo7802+Plwtcb6KsNA7WdziYDhm4byHOkLEI/svfw9inQWRJYNKyxczwZFwt8KHDUNZdcfH
dwiR9tDCH+c6x5kJdoeE/+WjK1N20PLU+LBZtcTSyYvFI0rr6yClIEwqwBu0B6lK3+93ww68e9LU
+ysHwmviZhPLRdL1Mor7qDR0oRFhUanchCifj1njf1Tp4ZXsWxTHT7rK+X1hO/OXKBhOpOFz1/nh
ZJ4EEYAlCTE/IafnX7G7nqW7P8U7VkrNQnNZuvOPnrwaYthbXIw0GgVoVON/9pQsJmTQrUX/zDuN
1XQiPMQAuKaNjJCbVc/ecuhorkSMOzD5FnLGL0NwZ6IRfqKKTtnrYTFhyx9h0jMEpZRywBCs3Dw9
ib0dGpqd3ciN1vGkwJ5ncARsTbix+K3c3AD71Tj7I6e+dBriJU2W/pqWUaVcOmgD/bskq1jNQgAI
BaH49H+uqVEqEKYZTLKMWuybBj4Ysl0eZmG14N1qlC/wLxayy2Xz1fvtBcx0K+mcxDf/Ou9tQjCi
3xf8mOWAXT2oJMQJ42XIGoTrwwYCMjDYVatOyQEuOUns0JyW2UQ6gpwcYsPNqOf8QWFJfUnzzI5e
Is6pPaib0hNARAQ5E9LgnsKntFvFwiro/8IyUbYnUrI24ZNdInisLnIqCn517Jwym+0WBr0+oVNu
5k8kXOZ+mBJwn12c+H/lj4iEfJGlmm+O39ElQs8CNgP3e2mUGn1mAo87A53LY3cAtH5tSUkch10O
uSXGokSNWv7ARfeeYEd5WCcIBpLV+2mxu31dDferlY0n3K139ZGiXwqYA4EfSAk9fLdTXgwOhVwl
ls8y2s72d2+STOKdkcPzjeMjlQ7Y1WO6qYZo/xYhi2x7e4V74MjVQ5fWfTZWbBUXvQngVOTgGK+f
puuIO10xD/O2OyFAT+dtjw8MSQZx/pm3fULE5cex5ZT0trEwi0UW+DLoEFSECRpWMjKeHrs2nJlG
mh8dw67sCkYg+Nx1UzQVfyxZDbErUuFjKfOpqBT6Tr1p/Y3Ub2DitxXdO/B8M8U9ZS9N/jh5WZ28
s/nI9uF4OkcgV9fiMF83AvCnAHRt7gRvs/IAoi3NNoAHqPXT9RJBNB/HEjAnenpHQpDU5uFDgasl
7X9xLQqj0ICFduiHbn1ylNmAJYqxeQKkx7lRmEHn58uOKQSg/td3zBHYeZzUSgzDmdKveLYLCn+8
tf53qnIV5VsJJkeqrFm+NTDGdp2zfL3PK/2GBM1tgVQgIFrP9f8njmf4muGNWjsCpJdG7Efgz13Q
YVzpzdyDRVs6OtJxlZr76cZmnEkL+gCW+4cka+MkuXbt80RLdtAh6/bKBWL5NJio3nFoLQPPrkZq
EHXEGYZOAs9NgQsSfb9G99VQNJD3tZQ3ZcG0+IJlqGu52Wprcu/Qndbj9yt+LVG6mOFi8zc61qRP
u+Fsx30ucRpU1TcZPryT5LSvI4LpYvO7fYWHJt3d90KhV+NxXfOhQq15hvErQpSs8fIsYinZDCjt
e7IY2I+uj34a+fxtvVOXWG+QnT8ihxYOIXDsBykpEEwsVKnjmTJGWeBfKHxQU06M9+aVe+o5WraK
0SBJGnT3BcXGxsPwwCKSx4o3PD8Zr4ZoMy8ConTOaJqOXJhjb55ruwf09V8EOv6MSEdZJ2UxbCid
aLMvMN9hl8odAL68KOSaOkt5IRrp+Axm8PbrRZhzHW8VamncGcBMFiTZ3MscsQc0NWgXenqB76gT
GYnUgyrc2bOegUVyIYxj+aOx0j8JzXo6IhzOivKxve0HAIGIh2/WjPUmbIZ/F+jFlk2isdzZtli1
mAd7xxDa4eeqcWnI7jfy+v+H5Td2vouUIf9tUpNb/kYnenpKm75i2SQNspdm4e27wMQWsYLA0oE6
imr8xiEnONiFQ7Msxqu5/r6aAbCH8dN5cdnpVFjZH97T6fAgTPzizWGDDMTJAG2rqLZwTmEvXIXu
Z1r45vDsDc1LiVDUzyGaeO8MViTUK2LgrihpfeF6hKxkm+WBv3Lp2hfs5MbO/XUaN2bxTA0cFEgI
tMK5iBDsaP/JY2uRCDjM7wDFi7xlRnBfYo8GhlQpLJ2AtFDwDY57bJlXUJrOE1CFTxSfSbeD4ju3
y8hWnnHIf6OJf85sN3zPMQULOF7yS/mZGZgXft0mVaLBLMgIlmqM9e5OKvVs6Q2GbrRKL8wYvJeR
f4qAuhRMdkZhNQ/69OXO8PQGcBewViHpyoW77uOQ3yS5gSfdLBFgPgy8nNcvwfEWYKDbRud3LRtl
QI+VWqKQIi0cgNERE7WyXkvBwP8bdzjF0l1goOhfFu+wsV5qLmxwLE3gTU3BCA3UsiyV0eRC/w8Z
EeKtqvlOn5nE4Jt8zrTDUbE5Aw2U0OpgCG9BKRBJVJ6YbsbnYFAX/XMQL8XrpTRXNN1FqSlDiyLm
yHeN7Ubbkhjj+M7qgq89/86Y9jymMwU7yjtmQaesrzvIMEuGUA7tP1gKLrovPBPVEVf3WP4jI4eD
LMTA+cQNvA/lZFTPipGiPjseb7ucAZ5+dSOGqXZ/rHWxFLLNUMOWVOQm9MsqjvbgeIvcl+Y2albx
XGMjIPM5Ej1/H+6JY4yYrgZzv95qi3usFBfmrxqRb50MCC2ESlxcdnVUIgg1oZ/jMP2NXkaTAU7i
jdAvctTvggKKuMtIZU/oHog9fSwCaU560K1LlKXp2Ji9rl1faUkOtjE2S5ZrJUbcgaB6+vwl6W+n
GbA+NMwupEPgPEeVIBhfL6peOLIsAbE4gMXFqqimgkwK04Aawrnw94VZl0lMgZnXzloZa4PkNXff
vuA9CmG7iDHb5Pvd4Mirw8dFmr2VQMWg0k3xIwGa+ulepy8GLFOqx5llLme4ZiXQbppzSJnS5/hG
tb9XlPRRtz2zOeMrFbI16p1n6Klhx+7zLzhR7/xdDeEXsHiOh9BAX18hP6fOmYO82BfZ6Vr6XAZP
j4y9heHR1Q7kMPtpgNhhuIxN3+OCn39hHsOZqG/mTgUeYDW4o8nJdUDAC9Qkv2TWBwsmaeZGpmbB
nt5a1yslUbyR7UVQpFWpaLrT3m3XWJ35Vnz35ywidRbx/E1zdCusvc75wE34cdDSoYOIjnsvWdkc
V+Lqfe02z09D3miU4h7sdDjNFGO+vCpUBNIVJ0bICtlzqksi+8eVEtvGstNRrl9LkMJ7i0RuJ0ye
WNc4g/tdsp5RRWKYezpslNb9idPCxzFcENq9EXBadjdbGaAGvNqFln5G7sYSl66M63Ub8k+il6w0
iLd0BE3KG0tnSFLIVCuPOW4svC4E8q4cTh3UBofwoBgvbIyCekLwBnXusYa7GWxFQYQFY9uJ72FA
Pvaw7YG30f7PH+t8t29F84CEyzjHOddP+tH/pN50UCqi0FZD7jaQoMBQuoAm/7nPFgK5L5MXh2JU
aWkKqdDWGKoYtDe+uhaTI/U5X71wGjynD5fO+LciAF9jw4LHBRvXA9QxewKCYB3b9F5SgGwSLwOM
dZyBUa26dWTCoJfxK+/wq3OvmNK4BqvBcTGVWjB/Uh3OjdCPDx/iEe1CK54/ODbASj9apbNarAhI
gmZ4qRhZFVIrm4K7BeuYFCwf4kUNz2O2j1lsewQK4kRy105UaNH7C9qlBnRD2ySpFbztJIJdbqTh
1g6mRbGdfWq8KvesaBv3/FPPmvtTFqhqM2s1JwNznVnjSqCnt2+fVM3PoD5q9qV2EFnsGhAWB06o
exUYe6vXPi6DVcp1tKv7O+2+OHyRDZpVDLnWMp/7mqJHXs0afqJ+/VtRnmEn7bb3m4KljXReREqt
mz5Cg5U8/3b/nbnryvLlx+Jy1ikvSePjHRW//P73r5Vo5uOMMgrzldsVZXSdLUgH4lw/+KhUgpeX
KNVjXsb5DkioH9UqSCmKit2iB7UXOZfjtKuqknz/nTVZrOKvpR9M96cv5z4ITTKI5VzWWRdc2uSS
/1r0zV6H+JAgV8Z4kmTq7EoEB2l9vzhb29Aavdw+XncfecTJ66q9+mRTSN+EeAC/8LAadfFtjMqw
aTanTmiabT2emQGyaXgPrgXAn6m8xGeSRY4aqmj6CgNpPe7zpSfFjV6rJxeCbG3NmPmg7HKYcsIv
7iW1WE27aVyPBMTnrauxH61avdifRr2knAXsVMpRPaGFTbumnko/FaZfU99yG4RQYU+E21oiQjHH
V/RStfjMKPTUihjFcdeOZNPx9qcsShKzAG4J8GHaomka2vJTxarYUaqkNc/HC7iKBIiAF/n7oxqL
wYN9WH2z9C1btHyknKcj1XWjZ0Fd+u0wP/xQrQmpIfaFjLYtc4a9otHHdIj4jazbX4hH4GZU8UMD
W3xSBR+rSsPF69M8Sty1aFWagn5DdijUH07Nz496cADXDTkj8WB8gSlX5qrF5kOnGd8ysXQxQ9kq
+FZuGoA7SdNP5L/o01PQ1Y67NNbnNWZMw0nqa340bvhqyVRgMXgEZ8HZhA7Z9AwA5Umf52VUjTGJ
G8NgDBVYjIijsgYu82QJAfqIelaSJMwlXEX4dX07itaCRwHSwdNj1Ldh1nCgD6LCveAgYyFOTPcN
cIgBPRbkByOyADnBLfOtJaZZFoBXGX2IsQdkGfKGTFl5rgIMET8PJYRMkfsp7o+eZo4FQDKwmZ1p
oFFqEhl4LD1XAuLcHQRnbw4mEqjOpBSP/ffRm9oJk66RqTgaZdSlN3O/qPCix0GTEaDaUmb54dLJ
lzZ6Qud5/Va/jw9xaQ/5Bwlt1bsHLdFUHLC3TMrQNotYS2G4pvQzOojYCc5/EPUdel1sYIyOR2hc
Fa9ZvRmvIFoYDfu5nLuWK4iLLIOL4PAxeQj3b8r2ema+hnYnRIs2rjeEeG7xC64SWSyo2IO1c7+J
cVAqt+8oYvGeMrhaMv4kaNTf7vOdpzlVc1rvN382ndc0pxqt6B2okdYkh0yk96ISp6NGPazt1cOZ
gf6/wB6A3di4BpQKmfwMpPtvP+zsNZJNfz74g3seTl7DTnlQCI5Dgxa86zSM9swL/fxC3ENj1wDF
3YveipHPTii5ok/WSi3Os9qQO3GRXAmhbYcV62EsSsuTarw1dQ8xmdQbzros56k0HBUZPq1lTUwJ
sWyu3XUd3LMISoNMqoiPWEEUe1UTVSjy+e+m/MlxsQf5Fh71R1GTMPLRDOWc42nP+Np+CX3DJcCm
W9BVEHOTTZyDN1HgHIgBMnTr+iO6R27qHvSdbV8yEMQYZBKFTROhdNsivX4+cRC8TdVx8ZNKHXTI
o+5bQdAZeIWHE+AvCzg/uK056H3kqSq10lTFeiYnn+S/REsjtt+x405DLngz0phK8kqbhoGT814B
6srYzgyrxhc3FxIwcHEAo2nHg+AHctiat2t4iXVkZoXINHNAn/Saxt5pGAiwiFIUaUSGkvrUsBKQ
+nsgGIGASYz4Iotfqb/R2hXpKQaBG/VP/GDhvZj19S+lhaGfFaxGX6vAlPRxD4IpmOisGrN3PDRC
/YG/kQGhUTKU8TZC5GoKhlJNJ2ln6RS+gR8SwOkUmmJKEDXbl7OVB8JCdZAtgnu93Wnj+5fE4TcA
J/inoHaQgtmx5X/jJs+4ZI2GS8Eo+RrWmwmAmk8cXMv6TFknsFNUAi7qAcraWq7F7uRbYvi0f19A
hUndj1u31qkuUUjQUGIprcY73qZGDWSQnXHIrquF3DQfl9/77eT4RstS7Y7ioUHqrxru4sLa/9j4
0rBT5d0y3U9qwnCLtLiK7+kzzzwvqs/l5scadfbK1T60e/fp+0jq5KTZLwtyEthOEYXWluTCQF/M
vDyaqshqndy4ZBh0qmJuRlK1ojDCqR4nZthhUcrs85rsQhDr8VVZgsxtmFIvBrUEV6gTeEqJDFH1
SU1rlI3ToLwbiJkw4wQIzMeQIdYVI5YLCSRVI+C+WE7e1OAfgPoAZe7q4ucjayCDvn+lDTbvxHNo
CdqwdWNfVX6UOzNX579DGqiiiCUDAqx7rfYSjUJfL3vYAy+/rhwIeEUPrPCTgIvM/qxt3YSVBhLd
kEpBjBRQNFuIn0+8LPuuV3v7ujnoZ6YRQZ5x9YVtIcHFec1+RyZErq899b/IwFiBTw9+0oiKRL4B
jDpvWVdtGPjV3+ZrbOUgy7qm7p7AeKnAPOQXpQCUNbuxw+Io/hAjzY4onEuWb9v608tPVecfVjS6
WCrTsEaQesmFXsdhrxy9iubcFudrwH+Uz4eZV8BPfP3/pDiENakhGhoHVT2TDtuj81+Di7qre5zQ
cXLK/vtN7lkKwM2TL9DUnTyS8OOKC7NhXo+7zEfyfFGSAg5STxEXgykadTEANgFQzirlSFM6G1i7
ID80HeIXpTl5Zlwm2kZiDDawpR6EssvgdIoC9cNxcyxy7cY2v5SZ+ybmE3Ds/u9JuwYdOslX95He
V6Hw4Pevh8Rx/TAtgCGE9IVbER0ON6MTdSHIAjsvH8lvOLgOf9RSLnoMFHM6scZ+uxcWDThYlMO9
KHAw2vDXtnUaQOcJBvrGHuFoPDJZRV03vbyQEbs0DpKH5Z/hmBHx2rrWQhs13goQMZwaWSqwAJaw
1LU1ITOQ446ItdIHXlIn6sttmTSkEc4w8aA/YvN2mZwWjx7e4igcHfSiCjW9v46KYUv3BbPhh7nU
ewyM8grwHEZn7tWi4vTJwz9LJhdiwUwDSB9ZNsjpVVhUaMEmJlezIfSNuBHrB13p8CuxpP6ZpD0r
fBp3iJYkw1JgaxMctwy6pOeun3l4fU4SnpWVtVq7tDVNfPhDHAfoDQ7fuS0Stt3TJHfwfj9YiOz8
Z31MbRldMKuoTWG6e8AEHtBaWDPu2HWRBmUjOosis3sTRhdkECntCvGJI3jOKvzjjbk5Vl9SQ1aV
K180SdkxJrVSI3PTG91n1wnoVo6/24A4NSobd2wEaQjt6gBFCWqeWmmCuxTOf2uAQpjTt7BNo8pW
x5XRWRolAYoohUT0FiEESN8vjS91Y/ta/C+YzV+KzJsJ6LEJmnUSHz4a/3j4s7oyDJZamU7lMGW3
2NZOrBLyxM5MirFt1Zqwd/LM0Ndw5lD+W1nDViRV3hlGYhLzmCmtymZkL+eNkw461bVpUnx+cVMq
YFzXRuLhrFrITAnEb9L8FGMi/vk2HVOqwxSn3QEwa110vH+tYCkVRHpsM4rSqqrsZuQFLdcXofnA
+9XXQp9+13GyWrsC4wqnrGeILdNN7Mg4S4D2/yTOfZI/KJkKEsciVHm8mCBDskQetiO5lgKEIBEP
Lw9EMWBnkmWXJ+aYvQm6lZusW5o4MCInRL8AQzFeTl72dOsPwY2+Kv/2+RJ0tlhxv7xdrwBMHAir
dDbvIxBhkqAqHTRJSmDbIJvD13n6Pb57kujbCENzoCFJOyofBcqaILjDORtAFOp/NRoYATEPsK6T
tqj9xAcfTyHcNfRx4tMD8pgLyG7i1521AQAmWonUw67oxQO69BObVC0owBdqYQenRdrkTcsArXoy
V/nI5cejunpqac///09sLhlpUrVbOZfhuik0509fVL4DlEOGtZOFtGZlEvCOBj7cia1X25oNIb8i
Mxh2clE0lroUJW67HS4AtbYJgPZQBqUDP97mau1YgkFKHPochkX1XSxXqYamUHjGspzIMqZ0qQsZ
qjttpx5DlFNzrVnv54glg3vnxGNzbL/KMOZk8MdRk4Dc78NN0uHrrklN4MLJ0E3ygbaFipIATAog
JLBwUYOxs/qRGXOgi8WVozy8QOb1qfDlXbWCTS1inSPvIloHWihvib/0Fbq+h50QxwGrv+1APAFS
7xt5AiCt+F/wgcwiDHsYZ7z7c0/YJE1RSYfnv3Ye3julvqb2TJac8YDqyWzdH9deOK2RY7dYlNjp
rRJF6jqPZOhBqstYPdAlGy7PywBxNa+sDfJAGJtNLwkLozXffMeqWhcOqzLNdu08hzzCo6fAb33u
gK5RayLMOtmlB8m87ECRYs4Hd/DMqz5iZqp6K5T3vldfyWCcwUTCWf6j0LWzlmdHtRyeG09FXtbd
6dhr5CGEjk3g3rJ7o0f43S931wCdwKklsfnKX3xTG/7t7pY8OmkWZvkz4am8PdHM0wB9eYTUOlVQ
t3myAOqE8bpUU+zSPgL9qdAWyjq7W5qmXQ4Mqu8WC1mgDToTjT+NkCb42o7x/qI9Up7INS5Ml727
B3WfA8I0F7u8NHwKMFV/PuQo0hpK8tavzAgTNHyMcGFVpzShzIdP6mnlu901bsF18F/VE31fPZGU
uXeFziOmVNTZvUWQNatPtNSTchCeUESf015gTgScUv/1pOXqn9ypn/nmojoM68UipgT2WzeREWV2
ankbbgvk0B03hSHoPBbvimEbNHpjkFPtUx891vH2E9Is9rraZCh7n4L2TEHo0zf2ruMoX2nMSL8w
7V/zZtLHr9yqSy30mYoQZBAu9oJhLUWDLhe16P0FIKCixaYX9x3Xf5MZ/WsCJ/k80ZblqesaGOsi
cspaOhfiB4umwbdhpFWp7qEOsFz/1gvj/fGkjyOVytAE3c3EWrahz3ENU9ob1Ltv47nT25O3x8Lk
bvmsK2To6F64uIHFq0+Jguf5GOhfMwUpAgpB8lTXsPW5gK5/3v4pOe8IDIfRfjh8s3PiGNJal/Xr
6IZSGdrkzu+I+Z5nL5e9u6N6tAfCKHMAg/9QGzFuRwmb4TYs8+mphTTDy1m/KCNhgrL+F79dgCsg
2oqMP+ctdpCImPn8nZJksnxqMkuguEdmny9Ox3PBytf+56dSRvxmyU+HtfO/UhxAha2DT0L2Fr5L
DdVO1w0F/BXgEb45YxDuU8Y1Jcu4crlJ+Yy1Eg/UfQll3xcbAECX6l6xKsINimlj6CtwbcoBqIGw
SneqP8wwlO5LmRsavTpTPDhr/08VUUTZhuERk2vNlPfWTTGfGBvVah2Uv8RfhqomMNPTIw461jtg
vsb6NX5NVUGCH4HyKCsdjaExC6mvcl9DplDRhMWhYkHtaNI2HFTQnJihD246baWddwu613tf0ukP
MKpNGA1BqWd87MC+BoLU+qFVhes/kNoAt/U+fXXfdJJBH/A/iCoKgn2FMAzpdRNg6gXGY7+MSSyF
653Z41zt3LUrHIa95PuyptvE2BHiLo0etSI83mNjMUP126WSeFJFBWFO8908Unb3XnL8nUzgOsce
mBeqQ/FTN8MIuB0pEZX7RTyqnnfDi3ik3xI8hkCHDdZWl8qPLjZYfZaQZIG8P6rQP/yMPMnvZ1sl
iL/uz4SQw4bLyxLpVRuitbm8os75b+lJZMq8UnlEkW4IZE2ebD3NwLgD2q6Gy0E+sSCg4hhPt5JL
huG5J3ZVuUzK8rGNy/K+qYvc+8icwA6OLYICPvhF/pG1TnLbgJtfWcB8N0qbpqQEwCSLwYkcQzsG
tk2Hm/RKQf8tZsJoA4fFGrlJQyXOACGach8Ujv8TZUwmWJIDieJAP+hwZapaqHO/VPUCutmJqXEs
S6iybHXZxR9OMLBnZVFyH6mXAkQflyOwbR9PtbzkwJNPPXNU7QEk/0I5E4Fx3ubHeCUe+p5TsdJl
6+nk9vCztRtZBnF1XKETpcE8lCf4mFzQavbGlL7R2+2Hb+jcDY4LVDpJmeuXw3B+If8DBW2L3tEh
MJsRgbGScDrZl02fvwsqiSQADSDf4vbqwB194ZyWcZS6levDRZ9Dr2dQH4hauQ2toe4T0EyG8Ve7
kJF0KLE4zOto+fOwGPWdUBKLBQLY+/MXz6sXmRj8aEVS6j+NS2djuOoPMs/hjIL90F6UmMMOj0d5
6vHRcTLdQiwZsnvFjIE64oIUp39zUqWuiNzHeIKnvO6QhcmbChug/c3Xn3jZWexjlVitbi3FQlBk
TiOGHqEmWDRCy6pFsV/9yVy7EsQjb00LdkgsdQjr6fTkZmH+o/ZKIINkFwpHDx/6A/iYLfAcRiWk
zTrVt25yLQ8zQCxjijxBVSNAg0sggZVDliWQBHkC6sWh2dI4J0PrIHmZZ++VabEO/HEi/wfyFyzp
yLz58+Lo+Hzoy6w9su5OiOkTfH40kh/IfhlT1vTf4eauUTnlqPKACzh2yokXdAh59TniCCm0YVjo
udImZ1xe5aJTTgpqpG30CM5cJxDxj+X1YdhfY3oAEjS0bgrwXXx5IrrAe5bfM6V0SW+aenNljHiJ
Wn7aKvI1HDJpMrh9sI3CuxLspUGzofH2EOUrrAudXfntprex++xYJgHoahr8TteHWAu8xL1/sVVE
tpr8NHNh84r9gnc+wMQ8FMHPqu2rRjUwznB/urjRwtIKih1i1rvY7UjNK1QnLEExcLItL9Vub+rK
+i1DniaPHYUz9ESVnwA9paDaojgWcqYUewXKDLoRNBhzkKqop4z3kHZgnxiTI+K5dD3GcWQ+kEN7
71VTkMuh1VuCjgKqBB3M5qxDdlfQhp+LPPYNFjWazduMALNmIi2xU08CdrUPV2TP57nPwUIR2dhs
Lplx8q8XlpPaHITqOh3+oW8b6a4ZvGHFncn8xqCrQmzShwW4yIRvs8tgNixlHn9QiCyvN6DBqdOu
r9XlZ1J74VOQ/NX0bgiE9ucBEgFsVE8F8+jQYzmTIg0uNvIT1hbAni7lHhHgDKLYvs0ODkR4FDwi
+w0kV1WajHeYkINtM6WQt/+Vgnb03Xd1W9BzVAXfStZSU+KWqemLobk9ZDKb62S4YeVVRrTMd79z
w083xAqXuVbH1sH3oiRGJmXqRo/jOvsQ3VIp19TN4HDsiCuGI7c1vo9R+fyc8C8hx6POFcgYZrd8
ES7KhxqiJhIJOP5GYr2P8xQTzd7IK31L1HpQnGMPvGohxObUvaoaQ8QIKO9SUw5cpuFfMcLfbmEs
4yfNlLglxjF+3v2+w2MBeLSqJnhP4p5EwGUqhcBsFunh2QoUpnIzz0vijV1+o+Uek7nCo7xpcujr
6jbEjrCd9NlggB63Lgr3Gp4vkhfL6Q7O9IQ2b9Tj249oyDLo2MUWsT7aPBShxXDWmjiMYGfiVmzj
Mt+ks/UIjmbOtKN1CD+LDNWpBJMaY48/2CHJULbQplKPuycvM0A9JTls1y48QNrlWBE0V6MPoCKM
dA+O0hmPT5UbKwz6Qcx+fiOIt4xOBgQFsoIY7UWHWu1r7J8LyYlVlkjIGblNpBNOnGfATeYltV8u
obV9xNsCbLWjPYlE3ixhnT3YuAeeXm4hPEr76vEBDZjtNQQfOHVRSrja1E+JPun92cHBVtJ8ZEx9
2ZbhLUN0bHcO1GsExN0J+4LFuniu8Hsu60Az53CjcCsRDxXTDGvO/aazuQNAP9Ec/4eEeBNgJcic
BO8gW04A3jnMaI9t2JKNmL38An4/Lze1oLEWH+2Qbri6xg75SsS7iSqqHdiGDqenOExiPw9mT2qP
1aEgBnPumSHVhVWAPqxVhmUFmRk19lFDOPWuvgp3PTTwpPJNQd9v+ICzbkizqiptrSNeGskhrWPB
aMJpyE34nyqJvezJgusNDJWr2JjuAyDTr4HZfWQcgyHr303L/6W3k0RweoxOBggXYgb/UQGaUOvt
DpMIZAxNZkyXPBD+4H4pleJzYcRZM+kvtMjXufxBoz3rq5a4h2kxx9zeNz04c3AdHGls5AmjPKL9
3bFMh4+vlpnllQyrrCQM7igSEVOKEfbfN80+kIo5U92lPcRZT47+BxbOvbAtxYxUws5uS8h+QPa7
oh6v5lusUqkr+qVgbXa/oN2+C4AdjIu1XZ4x9cx17sxhbd1rTtYoil7O2+B0Zt5UZOkeoDnBAUyP
kytyXDmoXWzB2YAGmYNHE8FiEi65oqMukQTJOSUJWZQ2NwISrgJ5Vjcnh2LNWkbkFysEZRXNeVxa
Onesd+pBVqW0zwA0cI90YpoBjSOJp2Yu4D9OHbJ0A1kjSGYSAnCtjZJOjscWpT7wT6NoiOtBmE89
4BTSLsJtchZ6Xyvp81f7ZFKot9ffO2glONYeQeB+o6m/0Gr51oihXw4uMlxLDLg06Mixh8RPfX7D
+qLA4+OQs3zXqqFgL+erhM7CcZOakBM5ZZuTkWHEgy1CNbf+iVenHVBIuKnu5OQlQmIs7rCXdYYC
oJHIZJndXawvrncCwqRnJlpEZ7xI0M4mBy4PdGqj3MXBKJKrH58Cx5124ovy75j8qaMso/NUwlCA
oY4WwMExjz2ZF++BgutFzfH/e7tzVJoerpYatIAR8+JDP8T0PlkTOI8ZFNvQzTByLss/xLY3kTVO
RYaTDthMa6YsOm2QQ77EUX6ySjW3pP3WQfMn358XQgLN/GVYEyB+L3NurbBEBnnIu2zMXOr7gukn
Q2GZRuAsXbK9sVH6tnIheSC2kZ/c3QVBVLdrXDzVt78Abi4m14gagTb2sIjAv1IRfxxNb2w+YqUG
QW2jF10A48/TaJEFgE8m/YHqRAxQ9xRP2oTbzB+8i8VbM1QsDb0eteZJpakkcVl5Hv1GMIk7Dq40
j9sL8PMFlBzSUP3RyTxXiCeYy9MSnNGqZj6d1VKGMp3ZTMN1bj2t5+sRREJFwTFhJ3K5AmebUmOu
yCoCOx4EOu98rel6/v3Yzp4Q7vnYf1jBzZvxNkIEkyYxYdcIlKFrsvs8rR9wTahuY9TXDjSYwPCw
fyBOO66+W/QLSZf+ulll065wJt0Six50qKrWJ+dKz0i+i13kK5EQFMVHkg76OE3sXMCe8ywzrgv+
rTQr/yOR00EaTljghFVqTZq9cCk+MiC/uIwKj8hjdpkZ8kB3zUEFbWJT2Gj28qB1FZgwRh6t2qPB
wciBGFjTZ+mjlXNnSSNa15tM/uK3Z1xIQnb5kd4TZCW93Hk1zaO1OofnMQJ8kSvo8fUDfvMfmFjn
LdPTPK2SuQTADKfdoG37pm/fSEDITsb4P8TfG3u78jAgeT1rjni5YPUi3HLMyyXmmuN7Hq6p2C2R
Ta7CiZG9xix2vM2hEl+IVPQznPe0+2z8VgN13BkyKXCRT2Tkcb/LZmtpH761GKl8ExTGFSVaAxeb
XA6FVzyp2ahTpsbQWqsIut4g1KN+fHp5QFtlAJrBU69j1dbjnDtEjs8Iff5WC2Rqvyt2rSlBrYfl
wbO3d/AZjFJVqu/E8k2TmZd+UpNmRca3Bxo8G6RY9Rd7GU50VkNZmwwPCAyW3zJX4SjPrL++jxvZ
+B7J2ivVcUx7h+bfAbJUCytTq4xFsBaKt8sO16sRvmxSmUFuySJrBsnul3MPkNNVYiT9vN32nSOy
6YIOOJPKOhyI3JhN9SjFa9/d0OOthfiP/VfbQxcUQK3pgnGb0l1p5UtPqEOI7W4Yc5APFqT0bOKe
pF/oXXhgkg+5OzPGsQm49rYxBJQvAXPofHQxLtdp3HV5IF5bGKzSgFZ84YSTDlcPoCyCQ+IodxVq
cc/Vj7eBOSOwyt8877DRlnOQdnWhVtDLUZf5rVwAz2QWMWGAGUBRnwCgwDtXymT9o10KH+LKQ6nE
egDhLfWsg1gtnSK8k86G7MhzRTIFUBIKgZKF5ieZnXcANeBN4Ml2/06zfo5cgps04heVRtoStHUl
D/C+OA7DRULYUohgj0JWRWt9Skv2D07Gw/TDkDKW8eQU+BI/THIMvijvrX7wE4iOgEx2b7AYAB6c
EWywQV+mJyuaOLSL1sFmy7BI6iH5pbEYWQmqMpXp8PGhV0u4vYDHvHsS6PlO6jVKR5kL/2mRr9T+
nXLgHpnUOCug+5gJb/bo72Nvh7zi9Qk5VgR2VXqIxaEYzYOppQz5kRk1dWbXFBrZBPVxT31P5zWh
ghQpGkAxF5L6mPZf25I3+n6+o2fE5DuH7EhKwEH+NADeKL/Dw4+ECsNkjFPnwzdhu9rgVI0A1OS+
jKsQG8aRyZRs/jqCKTZkOcWcbpRBMZ0zEA40a3+rlUThLrid6U2Gbnz9yFNkQOtTG/UWOaUpGDcM
F4Z/+VTInn5Z1pVb3rs4PYlaWU0s4ikNw2VscQzWvbfNHSpGgotYZBTLJ39JmneXQ6hMlY6YfPD0
ktyUOpboGmkwx0t4eaDx1Uke3mYsdIdkYxcBwm1KqVdkhiB2OglQ5HdvcJtCQdfRGV+lN6eR0xfl
BYIjA2eziLP9D/TowiKmZFl1npPVvMB7gbny01gG2UihtO0J4zU0QaGR5E8c034eVYzVqmUIISW7
eTjBfYpxVG55jtkJkCN0wmMtaQwKu7ff+K+8WzY85HeswEqqTfIzurYR28WzLppmKMAiWpTjbSca
JX7QS26or6alTyhihZxGzqeEu2vlqdkkc8i46b+EKVPDmLG9FDq54WOOvLPxPECmJvEmho6UCVWS
lXm5wL6X3khcMRxYIhJEifSnwlg9b6RDDIsZZgxmkJxGL7lndVsl7DKi3x/8bU5IGtvxct+zQwUi
WCIskbmJig11rTaalqPZKz7QpRT/fq6EZ8lY2cqx5wDHYWKXvNKdZEoYk6d18HE5onpQPSvZNj/t
0yFzglikCF/H4irHfPbfTujfo/hLFxmXUdzX6sLPv0Mjvea6oBe6BWR2SHjcqF5d/rkDA4Ojjcjd
i5tQ+rxN5bgRIpPN3Z7WTP3x72V7Cwj4PtEzfvvxckgu4JY8hsHOhvZO/iogo/F44jOgcRz/ZtjF
LXmE6PsUBiNRLB39EyWhtLmV+gG+J1EYfD0tjE0OnF92BAhIxavLHoBaIsmZYTKI3h7kDPdi8MHB
RLA9O/utjMx3egzgrFL5v6irLh4c9SIekOW3R45GLnHmkU77JVUviDKQ4TWxTQejfrh4c7/rakC3
hjjtXAOfrlS25HRZWOHP1VI6mfJ1/e25PpNiHIryQW645dPlBUZcnUsIBlZKZHeL7q8nyyGh9cHX
IdUz0lHJOIPjljXyXHGcQEebsTt6O/pxAMm5g15Udwg4epzis064yE9REX7PVgHYy+le5E7qx+ow
WerYFeAKTiCrtIvR7yHJdL0X+quindUDQwDOTXgRj+hP5dG+sbsgwgwLDGUlB+Rnwexm1SkMuqZ/
gta+Nu412SMozRWhbCfPhcY086DPfnMkVMHs7ZHSKDCQgUvAwWUvV3iIpmFJkrRFgFAV1rYxIV1C
urihToTGoTKxYMhz1khMlvo7YCHoX8Nn90swXljTtrGBVRDLYRWfNP9LIpl6lzIfKJlyGXkD2jAx
ze1Z5BURR8JXjLji3WIBFToUOsInkihNwlOrsn0Lwq9AyCUkttnQFr6VJHCN3igSK4bFCLenIoEK
ZxdWoltwj8ig7bK14r6E33Tz/adtyiEqqWmY8UR0CTMfCcdff0CLPX2nFSQiu8B7fRuODj+r1suq
LvRE4Oh9iyFeBJ6hKJY4BxxJK0frJ8WiLooNUyj1raHKY181PCoyIRhe8Gs7CCK9Mno+t7HRv3Jp
pxPnx+gGX6z47gZkYSwLMkXtRby1eGJC3Q4qrNDHI5XcIJmmeDjN2sKIX9/gwS5B0EkbMYA6rUTn
4yTRWh10MQ1GNg0+vqL4njWRukUfSw65dMPZXYc+CxW8ej8PEb7jZmaGRDoFpXsKLS3dCKkFo5AW
FEPNm2cE1HM2gWsMdqyXYFQg+3+YyS/vTzbKzDj+hEHTnOe4inhq6ZshV72Jq9s4JevB0IvKDrkL
YRJK2mAaKZNcXPgsHYc/Llenm7KhC0BsXzTJMLVR4wNNwBRAKgIqYWrG7plLOIvJAwjnugKZHfEZ
A+QrmvcF4+jbkT9MWnTtqDqbqLhEN2+tecyKU5xRbC6SHaPLaMrabCokRdnZ33+CiLH4b8nrySWZ
1hvGW6sp+YG0hyeeeZf0cWwH5OqfByFzrHdXBm6NOyPoTysYXiSB8DyJDZUwX5gBagUMcb/PGbci
QOJjXmMTPnth+Qy/5KYJLJFLTXkHXqRLndz2XRKN6QnMIQnnBPO3A5Yal+YvLY4tjXATYuRW9R/0
Rd/nhI5zfgyVN8XCRwAwQqGp3j9zgvybpozXp0hvFZdQsSYFyRBNZy5qMKU3+9wfhQmswfMEmgMt
hIX1ndcFVbneqoHaPSni2Km0+3in7iCyg63Lxl6G7OUESj+DZYY91OSdFubH6pQqsoUrY3effM7m
sTCgmavITKZppTtiGoMcsD7acAlqE2c0CDnEHA6KjuKPcTtlZUh3HGVq1kwJe3VzkiCm/VB5c/9x
YoDqw74LghKa9vu157WMf/eLTgaDFA1zL//dURhVm47Vp40TeIP23hqJdHzls9TOLv30/hdatNC4
BxEDFe27J/+vgFBh6gmmSGaWzVvWKUBp2DpNR6f2j2CHIsjzWQRiAO9Dj3Aon+OzWLXjcuUeHZwW
TjsltjkGmyyOeniYJ7P23D6FVfz8NoR2eVbjbfa4n8yBTXpshTMAm97yLisQ/JZnQVuCV5KFVvyX
vfhLGJPXLl3exmQ0CqbKbE/kCYaQEwT034YGvAm92G3/DbI+Bo/WTkOFibzsxZ+h0tVfPX3wuvg3
JXGQmL5CmcrdnlMNKZoqbvkJTv65xbFolk9mySyT7Q7McXJ5KQZbU4B9P4OZzYI2EcTzfQl+F53J
Eg3WFMYU2G+1Jdd7TK69aZ4PlvUxqJVzG7IRbvQ3guIlQxgLaCu7QRT14PIvCd8F096+QmL2k/mV
46f7sRPbzOBumtFona5Bq0elnI076f3t45BbZ57RbNhPCwK7QDnLgwsFRaBnBp5BzM1MnC9mGyRm
tAPEwXrx157UV7Yl5q6IJ6gaxu1mncsTTISpVNHHIgnsFsTBKpg/9SMZyJk8LXsHaaR8bCaczRij
/xK5rtnv24tqCle1F4rjJMYq9tcj1EwXFv2/Le9EJA3KOJOvkI9dwcAXws6YhgSVQph3d2OIkzXr
6LdKGEWMx/C2jisIyjH60LHtzpoqveg7xek6l3tmnjsLkSrCaXmlVDQKt+LRLlgATT1Goc7VIRCo
auhwRMqnO4LcTAO3qqvcOmdrJdOT9dlOoqcTs+IcvTuxM5LPhun4xud2b0itq/9WSORxmO4k222S
rdGoJsisKGjd4ZA1Pyk/oIWTcPycaAa1gR1h08AJH7R/o4sfC0c2gOVG/g6ohpLTImtpRsXacg9U
ZmiW8FxWkYULlqHrJ+2xLzKDx0RzbRkG3LwdRvoghnQtc6OLMLlsCD9menDKZ0OHSPxdw9RNHCm1
QHBDi3wAfuqaPTGgyXT9XWZmjjjQQvEMsspMdZdK9yO640YweMp1N8cuia3uCdH17tJt/z7Gw9gk
la0IM78HadsiayEmSPKCKUblZl/5stLNYKOs7pwN4Vkpf9q+7aOWZ2jc8VkBZNWcnuehSbVzY9ac
sHrPKbqGATJnqmKj0Y0hZG86fMJwiBHkvV9i8o8mtX1xkp/56DzI8hC/lY4XgFwWhpRBiVxE693u
dpSaOboN92GxIjDzuLk25A36kk4vx1Ry4I5W9G4I03zQugp3GTYyKcLs0ASw6PZ4UFg51HnfGTVt
1CeuXtJtjUBptng4c217VxrdDpMArfcd/x05TjK7+m/2/KnnT7l7gNpliCwe0r15F9iTPIVwJ3QU
Lv7aPPumGIZejhrIZBNSu13t2GPIoWgsZNKFvUs46Or6Vi+W7Riu3b6eX5Q72/5WRNnu7EoppEWg
FE3bJp1uwZYVCh+gMrwQbQ4kuQ81P09euMzE8a0Ai6fpmfMzOzJuI1cn01D3f8Ij/k7xFSlVzgFl
VQwZwlm1JU7KohpzdPQFQQBHUJtRZQiByw4JPzEwtBClwA7gsdJwmBl56cvavqZBaJlCmscI5sJr
Q22OOjiiNtv0Vv6pfi/wdse8nqJ8sYbZsNw3+tVevp/pQ9KFk8tsssxsYAh3m32vNLg8fd6hKc/E
DV65RTDpeCisX5y1QcjD2iBaOc//lsA5buBpw0/rL4JGC+MBp+08KlvDv6SEw4zKXamD6ikviIoK
+UnN4sVlMhNqIgIkgpF8C6w0OrxU2//JPCmxaAgllNSwdcqRkTq2Lfs79TWpwWTq/SERT9vsiQ6q
rpWAluL/vQLbNJfM/JXSVHEy44X60kypVyxwsD7+SzpOhguTLgQP3sKjt9iumYGZDlUoVUebWMs/
paYHbls9pIvWCPu9rOCDKu4Qi9NToNrginxEfjT50Bknip84i28StxFi3++r6bSWt0hF62ZZKHc5
KtwzgOROiqTBG1zpCZOoNUNFbY4EozJBhnkIBfh5aPmVaxmQrhsYKo3hnharc5UUEgQH144Hr/K3
HmxDbELAro4IB5fcxXjWn1VuWCjFka84aLVLSbBFsC58h/PRDlTRSKPLq4YOSd39IQ4L7FX2mgKh
xpjnHWcLCsVB9XUELXE+ymNBFBtjkr6lbkTIU9OqOG+illl7cyImkD8Yszlkux48oT6JKE1DW6EK
ChOL4DWydDSSGnb5GZrREpICFJdJ8/xunF1DnzOJ3QkgdhNlnTXiiMHnabVKINElFT5aLgZ3if8a
lMP02Y4QVATFYx2/LdRaANYxNzYVM+nEZ9hz9OIoDqz6e1LdU0u7DaCEMrNH0ETaH8aKe1EALP4r
32dXTqYxP9LrHr0nZQifQS5d/rM3TLhg3p4VY5l9Xz34nZYAXBlp5lN3jZmYVaJ4LZTGIfc6b7Qc
a0DwamxI9ASRhf9L/0wk22EGu+R4/2rEvGNi8SWTHdKkJQA+DjF25zmCBPFbQZ9/UrOimYyt193/
eZlc1GGOVRv/kJdbDyvEOIvivkVmOntsurI1WjubF4NH8PXGmJJecFniOu1qbDPO+EvDzXShr7gY
7KHubfQFIJb7fmhheKQFONpNGhNg0SukuqXIJ6R2PM1k/AG94+xrNZQJcJ9gMfCuYJnK21hBOKvk
ZR9lT6TiInjrF6eYLxnIVuKZu4/WY4b1Q8EjuTI2cHC87VlYvisTYPFt2hXog1aI+BUalF02uzIR
174s+z+BWfMfRF2YDMaChV2h+O99RMxQebB6RrFkfY3aAdl164faVzqq5+I9BO1L6c12BplGLHYM
scg6Xy5v0nRC11+bVKJ4vfoGqh0nrdKY/I7kddc1wn1TelJoC1eKQI5MShDlFWXDI0gRL9tNFQSH
SkHbqmYSg4x2thXFoIc3ARvo6h+wFN4L+agyUgWVq+V/5HV2BxqypFt4+6znQQsr0mA5nGRyU7la
gH4PLJkA1F4do8T/ykez796EYrWN+L0yUgzXlIupUxadg8rPML+NG/qGhclr9JjB8oxKhhVjl1aK
Tza70nhe9gPdvsrg3jFoBHXrY03U34YwVZfQIpZQj2xpA560CXmnkadK7iY1OIbmxZkoWY7q19MV
te5omF+MQC9p1qsRI+x4/lt0GNnLzLoGalNCh1aRAVw+CJ3rkAkXxv2yCUyMstj47EJxkfjCWe9w
S7Nk/bT78kSic+4vGYrS2uPl26Y9Mz6GSY7OiSP4IVBcF8mfbPT2g5UO2CsGA6FjGv+vGU1fsAqs
Mji6Ji+0/RrSsm7KhhkhQUAycHhUzGnFUOLanddVQMhWXuMcEULOoTaJszNVbeQWJommSlEVAjN2
wjFXywRkEHy2Ck5XvKCRdxIVbBFgkjaEdpduX/VznmO1ePpYqFlMalCE1fbTuYG9Utma2U9A3Cbd
TotvjF9CU9sImhjPbE8Wyd9V+Fo6/LVnR9a+JzWUgRRMeNteCBqLLaovfgQt+ADumjO40VJP+Nqy
2XEhc+lncbVsMsRKIdOXU0tCaUEO884LYGoPh47VpbVeZAZSiRpeAjfIlZ0QDh40VAqwMJXMfZju
JLVT7ZrhUNRwH+hvfmZ6OzXD03kDlPd8i+sXM+T4VjdqyV0CPsJLJ8I8zJY2x9x/AT25YuLKv8Ug
VQY5tf5d9Svt2/zl+5oqbrNxeg2bxhfJJvPmbw/06SDcU+cDkmxQALZN7vNzJzfz+2DrlqZj6CjS
4doi+lBTINVnvxNJ0uV87yuG7S5e9h5mSmPgWIzVNJYmmKOUhUMY9XHHZZP8wTfsmWUo/SLoGd99
V5cMms01o7kndPNrSxSkJR6mXxP4icMOhSdLZ8me2+UmYmrNkx5a0yTcORvVIDFXDBv/GKuK4PIL
NxAyBeWD6zCZoJCTCfu7K+I55/wxtLxpMmi5HLXlnsEC0xlSWZmxn7maooFB84L2twOfBXryVihh
ZoU3OwVRxVLPp1OoxPHzNbww7ZIvwC6l+j5bZax7LzAy/WCzq/zSbefKfCL8jLRJpqJPbeomxXkP
JywELDCpWJEm808JUwT3hAZ8e/pVxGj3RT0ZZ09LxTIUFjcRaBbZjE7ax+A8lS3GgEbTmwjWhxeE
BRUgPagHsjob95TnNWcJR0x+p4HWYelGgB90CGfx7wBRw4w3jjXN3iqBHeM6H7QyEMBjk0Q2O9+t
G/0giRY2IageVWeG6O70IVllQSRvu1DBYu3QbwL7LKbZAAXL8k96yCQOFkFe0XsZ35e54gY1NIgC
NaTGmwnZ0QHL4VH4TSDB+8TSBmk2uvji6oWg50fCUiuf6xdPM5q9agpsh3/sf1+txQpf7ajMVhKS
St2Cj98w42/RmEtvF2h8QTlt1xgh0RgYcK/3DO7o2jAjW7O8P53PlThpWjdCefY1ep6ByGQHchLU
N5DAeE9xzMO1OhVCpM5I6M9QssNNIoCo/pWoSZvaGpIjFfJh3R8MlOKdcX43i7PWFjfwFgE1LW9e
sTcLc4BGIIhO7a/TQKH8ml4EHNkn8R4d0mXuPgkQ3lCBiO6DkQdIg5zDd9uBIBJTq7tCwm7LKroX
CnLQ7LuzM6BZKBrOYZjBvubUhlX+MhvSaCG9AmeyFxWKy71RZmnJlJkJY6iNJ9m7GoJagalaBF3a
4q78MCTgXZav1mIFxHDxGRYjz5rCz9Nu2KV879cS6V/0xrzsh3lJ8zFofy/+7qdiAc9PFWg6w06e
GyksnHon78+fdN+/CgcXhkqjsLn6dq/CWVga852zJF3jm0UIQWaD8YE6uJb5FOmBfWQnjNSUdqlZ
pxwvvcZxizo33rJoxE73l0jt3zU6Spxb1G2mP0NvDb8PCsqm3It2ugqd1MMv/hIftOQ02uZFom4p
GAHLG88sBle40wN+QFf/nVZ0ybpF7iPtyYmTVp4uAbYse7+PtRn9DmQwwlgBKtxsYMIWSP7Dx+zC
f33xfErmGYlPBSpghofOdi1dN18huXidOQDDU/jvwyxuCVhmEjZ+Fu+YQVK1/tdYtrKxAJoqBlz0
UJKDtGtxtWj69nWjJo4wMqEiAwzKlkXNiwlNfT3F9xAVRofGsq7Dy8Uom63ilVu6tE4ZJyHMVIlS
+crLEifYtdGEJuAGVOFqE0d5NRfKSMpQwBQsQWCj9KYQ4ykRJ13SAzIzwpZPlh9sWOQ9+lM/iM7N
ypJ3qgyBz8iM0YMWyBlfXI9VX9TOKlPwVvzVHBURCzGwLlz9BiKbfxb7BaGr/XDA1r0WycJyf783
DwAXMQ1+0kb7kO16JVYl2qLEg4xBAl3SIyBRwxpgLhEctPYzIc9V9AZ3ytN/5GX2oYsrOL+Vi1K3
DSr90nC5sEyRrNT1sGMXSvfRSv6UYK9SGL2If3iZGNU48uhbLvzOzNNfKu+B4XrVXtw9JG0PJZpE
yb6muGmGEd0VqBYfJKrasl3elr0J4KQ81b8IsgD20c9BvAzFbmRBfZqrgaoOEZBmhckWY+ZMBMJL
qiCnSIzSR3+FjSnwZ2S28p4ZbbagLQGEB7LdfLv5iCCmAmEE4FZgg9aCweXMf8fe0g9dg8P4Ykal
TWEtPrAXZ5+xrmeYnwmknl7WydMcVoXPrbzZPb95Y6RgSjgseRwId+zlbbFJFTh+xN/pQ+BrD1qQ
jQ2v8EulnSSAceaFbeafj+U8IUEyDkK49u7VjpygIQVtUeyUcxrvonR8wM5xmbuGkCFfD1Yb+OKC
cGqXA94hg55wHrtM/VyVmrRrzl/4gK5XCzfBw2vpUvd6mdnKESSmZJ23mhUmbI4SWrmKDWlnahrL
W5nvrlexQYef0ffAfXLaeParTppVupxhugpIhB6j/NJxe7OLfWwJgRtaPPWvDCdLFTDfrITqAKW+
KzRhJBbnOv7wvJ7rCWWx/cYET3tpagc/tkSD6Atge9C/EqezUZRFD8cT0CUiRqG/ARkIGyruRsW1
YGWwhr86cMWixQ/h+1BrZ9boF0tUFCQ4qqrTH9/TcK3mJ8xBpyyQp46HEtwzbMhKr/GZq6JO3gDD
2xmcmcGdkLkiD5GPHe4ROC2cafn/xeDWON0MI3sqU3ioZAuW0rAg7g1r7K4rT+zWMCEVh8XaFBES
aqz6iBoKPfjTTp40jakjUYOMEFcDVS4rBb07gEwopGTKwcKoNCMRHmC0VkdmbMI6I6uZwl2cN7ZQ
ug3FCjJMjEjTHbox2Kc96ha9wGIHJK6rFuHhPjEPzmq1PT54fPkciDBfoSdxizNjJFCI0KEU5r3u
AslA+ZnE+ArnhJRooRv+zl6BbqowImyw0FizfY4DbS6aGrOuxRH6nObcf9BQVWdgNltt8QVdH9bV
ZI2sJOxA/9vIlgxer55TUsQKEZ6gFSCmVw7FQZJNOmvg5eg240bZ3KIXmjgMJzuCJhlpW3ALgfKH
WAtq8v77xOmrGOGp2mLAkUFXjlJEXux9uXcHq0MSuZ4AuyOqEwID65Kw1TkNZwM65rQXe4yUbK2y
LP/cs0XEiQpQw8boCIq7VPerdKxKH+faODCbntHbgtsJJC6F0wKCn/UEZq5xYDmWg++yWG7LjBXX
BePpBPjBMGgl7eHqxhNvjRK3Uv74nVRt1mIIK71N6QR9BkVNkry6EsZvJ1vLQRkK6LHcn1/xeAVf
yX/1hfpgNGy6mPRu1BOP5qHU1NoEaHHTkocos43kc9RVIoUjwIyITwpTZTBHfIOBX6SJLV8rombu
GeHGKDxAhoS1RxovLDx/6aqgnn+WZ276FWMGKOerqCFUcEAt7oMmuhXp7/hFGVhufqzVok5U+taP
HD6TMn7Omwzir0KiRJFTN0yzN/bfWqYJS5jFYS+3uQCaIf9wdmWbkNOSkxCx9ljhFzzlD/7nfWVy
snOR1Ew4JMIVqtdXfTB2gOv4i+HnVDFcKU+k1b9hPRzUgkbL0ypgkM28gR2IEpbeVYSrZ51GYzB8
aUwH8Gi4chL+Gpe0FAIUO62w45xgpl7dIvMMk9gIXUCf+U94tE4QVbD+OPp5A0fD7Ok4xChTnKwE
r3kSX4GH9NyavY+f8yP/HSBSOjx7eNCV16Exru0i5jozHusW/byA6wPpkvyIT2vvnaCh2Ke8GrfK
1AA0lE87a2HYIb/T/URmiCaocHiY0H+v6/bo8eCNBDejFYmCnJ8sdaVUb9QbvXLt/nDW4KVpcLIa
6AwpQMxBLAY0TIwA/pMm610u6iNPW9dpNY/ecbPKhE/L05cpt6GmSWUHBWJP+vqiMTKPu2sfX6LH
uG4Jx10naB9eXE+WlBc9tbw8gHof71gcKM7yPVET3ORY+b7xUE9+jv65q1ZvXYQV29542TzW3sGW
amxamx/nVVpnfYKEe0Dczproaw4PO/RZkf9Lszpi3cam35JoA8+PGm4w4bHyr/6f/G+kVj3Fk37f
X3VAOa1Szp5mvZBwNBR3iYD1NwfrKokvQxbB254zo6IazPdPpZAE6v/DgM0qxF1AlSeZS0I1g/YS
jIYu0FRfsOYxN7TZVQjUWxxLq/1IjpcrWIKq462lilicdsf6LbF9vfNEVphL2QZdjRM/l3jpUvAA
ByNiol7H6UMSCa+oN3cR3VWwb1biYK+A56T8WfL9L8F7xMBM2xM5/pbvuM07NLa7e70zckkBQAXD
qeTmn+V7zh5M5lrAPSKZSb+9KuQD8Jwp2EqqM+tXpglhuya5y4aUvWHoZRhWJxSrAFeXDOqWQo+u
6D0uiNR7j4+jvhO2eu7EfjnvGutH6BXwEAT4eC/zkU1N6eisOAq2Y1Sr+4m2eGDlvrK2L8ztu5CV
X0usrgDc3L/rrXpPPvBtXyETbfkcX8JSdysBjoVuFf1IeH7pZIAq4DkqwTm6b8issCf6WsISod/k
RoxqtO5nlyv1HLEpJffJ1OOb1+kY6t3Ajk7sqW6MAurdW9/ctiqlr5uC/GjO5SyLtVhH7wO59jCM
tcoIsLPmtDLTOf6pC9ovSisQvfc5739RM01BjZY1qaZx/xJ4S5cT2d7RVEt8yYsmJ2LNTEvql2jB
OQi8AmoGvxgvCATWNnypYsip7czuI27RRz4dRRW3tp6Hf7jrbUz51wdkfPRm5/hMDqTef35JtxgI
28EFpMi1QNZ03rGaGB08RjgifTkQyfxkUDX/Q4FY1uDbvb0BjGBL1kj21LPYToZb3MyJ39eV4ToT
iqnZTE0r8LY81AhDxEB9h/nJz2JqPeYTInTEAzWiH7xoen79QpmgXtNTuPDHl9eSEOxYvhvnOi2D
2V2tNIpmkPO5VkoRjCuUtYtI0N5KU3DQaLZhhdEQkV7OIlUMH4CF1WLAkOj5ksZkWw2OdEuYg34Y
jz7klc0Md+ICbMvNUuO2wSZ47Z4fw/Hz8qP9UiE+e6yG8+pjlRmIrxe3X47HekfhrYjAOx/cH+LC
UXpDH4MS9st76WpySs2L6f46zCnjxsB3bGbVjiu/isgLs9bXkyh6BwXlCTEbTq3GmqLUQQ/R7wZ/
HSxJOmOlIFOSZrcmxH2XMqt2Ie+Iz82UHG/2XswIarBthc3yXge67o038keW8bBTS/zuEJL7K5jx
N8yz6IzuDt68i/o6eUtUgkHIMnzSW66KSZ8lCniJ4MsAwT2QvoWMoxhaaplCZiAGMdC+QUyDdF31
4mlej336mjTOM4HYnIVLmJ/GFmkO97ygV4ueWUB/3a6hX8uf/sEr2ZiKtp+PQKLWU3Y9mVt0Eieu
7NIBn+EIPtmhGgiVOeQJ5ST4b53gJrC9QawSywhtrg7oXtff5VHCC5/pjAumWRyIUQxKlOZEPbhj
7XDO0CI+gatnm4byptLIiXmXyc49vxKW6MNgWRjSzjPLF3yHJ4Bgc6RZhhrG8uRnR0zFAHG142il
yKZoEO9d/8kV3EbUTUGlsnC3f2j/3mr6MtLEbRFrjoIHQCiRS9K2qCSO18ULAersLD3pzsfdsSQL
nMYE9m2yKUyuxAvfr7STLAcTTQY2pI8cdoRU5umJOMCZ6OHRuBfS3nssX1F9aHDJ+bleAo8hxKF1
9u/C17m979gjcVLfsX83qbVGKCrO3tmcRnDLexwxkVUcjpFPA+kE2W9QUINiOlQ5GzFgY7E2Azwl
+4to4kPt/v7KYJLezlMsCqA5Pj5mMbuMFaqxXeq2NchANdc1+reb2fzMUdAJn47XOHXU88vC+GSi
eaovUzKMkurUzpSrPD99Tc/kk9cEDjjpzRE+ielNHQWBUwPwY1AgLmvqm94LW8OjGIZgSAN323ZL
dR720qXXgSo8Iew06zKMuv1uayX+kSdrAaY+1OkHRQ5nfeGNNKUFFxB69NTzn+0PdNriqx2cZqfg
dReeaoKytUKAtyy1v8MHbLKXCiPndWbDWPvTsH95Z/bASVCnY9L2cqkM1e+T9ILINlJT6N6dfulo
V0JN6KetcaSFknlOTxByO40Qf3leunnr3Nz0YDIxOMdNHlXqj74G7xxyAH+rRh4bLn536K1q8TrS
Un0w3Kaldg7jOzTqUffi6B2krpVEi/LVPHdKPgFmqGJcziCt1TcfbVZ5xgqJKfgD7AKrzzpgWBL3
UHbth4ezBy++sDpKW1Qj/vg6PH3TrK5OLu+EOm3K9IVS5aWkXL/nR5zrRGdlnBwDh0jbCHChjFmE
tZBxSHafx7iCNdtMFVO3c5nCQQLukkBTQ9TndX5nHkhSnOkt7wBoOO5oAWaF0dq69fwyacsEP5dp
aqTIoud07B+Es2BWFegZZ4boY97UQ0YOfUGNyes16VlSmKjaQ9FNmlv/2UXsPdqwj89mEhPU+a21
DFbncPOUhFKMpr4JjLnWJFojsaRpB3Oxcyuo3MYrjC/2+q1UB7baSQfB4MJCqT4VgIVrgO6BSKkT
/gXXoXTA2GLJHNJtIgnR7b1yLyXW9xSHsT5B84IefzatynAdSBwNoxAoFXF4v9WWAI29s+ii/nE1
H84QuqXwvjRV3/EHjakYzU122IqbI3U2z/a2dVORsHFlPYZFoaf0su/ndwHv+rss8rvxzJDQyCEk
KKY+lT2ap3JIuCiudhp4WGggQ9RZSlbrlQ1cfHmcU9o//drA6kQucvtYftCXQxkVqf/rXQZuMsKm
2HMMkjOn6CDqkvyT0dfJRxgP4eoU5eYsidUVyLjbXx2uMr0x43NAbfsTD3EmXOF8vlKshrJjQRqz
AHHD4r7PAWgC4licv7pgXEGCxexUESVu1vL7q8UpZn4EeeooO7yw+yj5ZDAUywknDuscFI0NnZFu
eZPVBJreR2nFdVVGzBtBX+f37R/KxHHtipyGqpbRKomI1/wo++ejCMwntdb2n4+si53hvIq/De/W
DkxIcTVcS2Ri+KOAn23Y/oa/K+iYq9WaKLQOMuUh0gaMfMdxLCsPv7FJ/mL+AjyOdXvFD7g9SjSL
Ql3XKwGlP0azFiE+i349rUFCB0ui+SsiYv2txr8n3KL8T7GKLy0IJLC8oVPg1GYCRQdlIKuoaEP5
WxZTAf8kKKTFPU6Eq+haX/YJKixoRWqISkGo7ptlkHzN0SXvUSJ2hWjBV5O0xBRgKJ1VKHq3sx8F
62X523l8AzGX2FFbqoMuiY00L8LfaMODjlpZ85efyED5Y2WkUt7/+hmHXLLJEWgr2nmQvMIyYgSm
5GpdxUrMQWwaw30kl/ST37eVUs2ICAX1QvImGoqRoKXQGqXLeJbOdboIyMI3f/2xvMnMWcbwzL0F
Sf+HU4Ixl2hisTibBXCdG4PGEQYMer9pM+IzRTX5oBB0O0Omf5Te2abbbis7k5ssIAEOy4MUrKtM
ktdNM9zSQo2HuEBCwsWyRIAZbyA6m77j9tsztf5IzwNpbEc/fXYbmrlgC4q80siWONlhTtMq1Yi7
paTnSgEjra6AwUtofkT0TekkPYtcX806sU+TyUF6iKnkP9LP2TgBkKWYfDTCd15Qg0wl21j+qsNL
dTICUiHBgNBTXHO/0uwGW0++h0PKnpNEjFLyeHNsAQtWNGXFuPGj8Qy+8gWtix3tVG7PpgFj+Jl5
4HzRmejMc+I0ektn3hbPpxW8ntLKq4EIZyMTOdtp+NnQyvfSOLvZ7+8TXRsRxKRHE7Xa7HpBug1e
UxtLrAQxNthXgN5vPUQZ78UIO/RRGxA12Qc8UrjKGy+dW505Njgf/g4aGZRpo3wkmYT8siUj+C3k
hYeGOgHwKRHdhuefOh1AePKls25EP/LyW9DvzDCQ5JAX6cjoupj+2d+rbx9LNmsNytl4DdTAJgFm
kl4yqqDAl3yn2x8/BWZ8vXYtgskZmZ0p/dJjW/RSjJK13SW674LfplC9S3SwuoYVPmBhctC0TIes
yhtA5CVw1GTiHzkb2/Xsp0OCKV45tfYklqW/HDYjypXOhInYpj25T4SnKTeRLY/zj+QHvT4M2qzL
ED1Pzs4UCncemI2cN0EBmZuDgaI5MWeQs9UWvJLL41m86b7m7tVeQxPhuVVSbC1e6CZFRudR8Ftw
DD5cVrwXEJxTcOL29nYTgAlKdecjmjNlFiun4oVDTaJ8qakkHKEO2lh+8N4IHLfOVkfoDTDH54ui
YChYP4X9PQy8ECVYjMiJK99EdU41a5fcehmcnpqkT/EH6vKaKCghF/2xpaS93eTWGkEf4DRw8Bcn
K0CfE1r8Tnbma+GELIMBKiH/T3Sie7yq0h6kZ1Qq59c9FXeLQEfg8S6QRoOU7kvd3qEdmHsG9REF
4BueuRXW+h+S5UmopQbP3x8UjYhKxBQw7+7svu2cQKINSrUbdOKUSO4z7paIOcRb135XeaSdM6Ax
2Dg5ZGJ/IVjncKK6R5q92k6IM1Dns4E4aYV0NCHyAYQYMe3ZML0h6hSydWXOd9RUDqo5sg3zd6N8
wS5gbn+qW6fV4+Pk2sIawiapop4/MDz6pfeKKOuq4HhipHV633/6EaDJ9CAiVHAz3n+B7/xwEfFi
RtIWyrB09mBIGrlSft36zp0pG6lDG31aNNu68qHf5pDfvoyDVqhdwkzCEbexyA/3BISCLFTeMbOt
IVAXwHBn3PZcWIIApNy3Bx2v72ejdjhCtL6sx7sonXHhxcgtlx5SCwdIR/jXZeQbD0vL/heeNz5w
iKz6uvadgPw60FjfREDKB/0BLg4nZ8C+9YXor5s3cUTrT+vLo6AkRob4R4yKDynyombA17ovc8H4
YqmxpyGRlgTouyrVxzwMcb5bHDkEHH5nAUF1sZ79tv7LsgMvfgsJ+yd660Jmyuewk+n9Hh+j0K48
GeDq19zCkhfGLijo7r9PB4txtc7g3eYacKM9QdkJ2fEVJtcBzykTQEjjyKiv7mOoULfYUZ+B4iTb
dry36TXo6RCFE7ERpHGvSX0nZqPdRc/F+Aek541iHmEkUUtTLhw6A1WOTniCUdqKEzhgaAucCNiW
9GVZk/IoKpIncH48NXv9BBVJWBVi1x/+Iajzhw14BL79azWTcMEfEq8MKO7zIe2QsPzC09jpcPf9
vGf/WNLvNhGj1fbfNkm9mW/cCfU7OE3Y+15oVwr5OREwIAAKJZn2V6/6iTbXtANxvZEK6LFA43w3
JHq4NkckGUAIdLAQ5bw0L2hiZ7Q5QuBj6tDJDc9SSwM40YeLFJm6QV6uxoiCZDO7tNofHsQRZQpI
YLX6PVfOOWqyh8nvT2ETyTYnYPY8B7t2uzKDKurnnafBQGv5dc2JKffm4xIUxMykyJWSWXGGvSkT
w0GPQ7+pZbwtikXL8reD/9AtNYaWjsmZ8/PNLEXbKRLYK0vPYFu6oPGt7J72Jg2Jkv4cG+8Nmp+8
raCwLMw1Cht30ZVKZ5NUpLtz88wMDZv4ocVUuYWRSSMNrMbeFIahVzeL5s+kwApGv/Lcwmbj+S/C
uz8NiAueySZ+hBZCp8mamsI6OGzFpUSjPBndENekJPDuZsHkwuxE5Fl+31Ks9KE+ufCnQC/YCBCN
4tvlb8LcQmMyQDhdLaIxCQx8OAIx1q92oudDTKCoOkJoSph1vMJGlgZE1fwYshFOrnfau7c0xkWc
VUHKgW1HQcxrFG0Dz7+DhGeFaubfQPinkGBUWcXPHBjFo5oWILJ6PzfRwMQZE+7ZIfJ3X7vFGsuA
qxIHWuMnjXcCskkA91J5luhiekDSQjpY15WqNiKhlS3rSHlsWqYIrhFs6N8TqugjK4KTTUqZqu1R
IY680C6RmqmwNserKm0WDp0mfgBoyoHmX7qG5wU5Lf6oVzFoCJKAjO2zifH6PYlIJpBibyLegAJd
TYODdyuvSwVPdhXU5/8tIAiUgy+stnjwuQRn2kdDPPz3X+dz/WVEMwzupLdrUQ/PVRFM2q9XcVht
EMHZF1EFSfM7bPj7eyDZyuKebk+gxkt0m5xYZLfbOEwlBI+klxqxLNi21zgfhpBRuwatErl+/4n7
4bdho0bx2+VIE/f9jqrU9gc6fxRt7uiy/gQhrgkAO0vRvxmptoz0E8K8bgOyrlohGvt04HrhuILZ
P1mYcvcSU9Ixo5i8o/hte7AKimGkCGpU4VnFj7qxt/t3zNJ+qQVX7Xo5y+4zj8960rTesSMcaSEH
c1ytV4VpXGnA96deG0esRxgmQek4YWB9vFDsmwhEQlTruPdlNcNPbg1ft4jhutyHTk3ftiHQ9jt7
8+RiR1WJd/qlgLw0aUzWkivZRsb3uDYFKq/Y0lIepKvMS0flXwNJPYwdEten5DrRDO78cVU86ATz
S3+ecVOmeUwpG68nopPlTJM2d4/SSXniVHf1zK8jLJORbYcirCQJnvtN3OXnbazglgu8GR6cIUV5
Fxtl+yHNz38S8cxp7zWpxa7DKk1Oc0orxylfK50cZjiEDzhVYJAnakBUDyo9385SXr2+nOMdEFAI
q784b+TZwtD+EqdDHzFUAYqJcBIf8uFJ2t793OMW9G26lsZH4BNnFIpS0eyzgPpQrCsewvyfIOJG
eKYC8EvTY5qqH8G0qygfBZas5m5FbMyUdytG1959aOFsvqLn0hNYxBWPzI5dmDlvsvVwl5JflbAG
AbObx5AdqCPeCMYYHbvjoJHHpWvP8wMEiXH9hrG1qPZsELd7lJRhLtDFSriUX6rM6YCer6rGLN19
7z6E2bxbaGmo+h+4AQT3AG01XkyJoEi+SkR7nSU20nQA52OWGu+3iiKOd2F03sVYEWLPwSzCC0Tx
EHJQn27IuTBsDQlhKrakBg1O/PnxFesHIVC4mMNFpIb0JryIhZAIaTBMb6KeEep6DhcM5RWqM6Ng
1eaf0yE15pkytONs2ixfeEflzQ8HV8D8c3Yy+3h1HdBNiN2ESNWbKxuhJceelPGfDjVYoC4TnA/0
ueUak0TV3G3/HgRzrcckKDk18+m8mccsWpLisEDDcOqzKcFrwC7QaCsOjmbgZ92QbeNwtRuT0cdo
pwPdhfnQUD2kDV3wxXdlN0ENZNOZHeAFSkyGa7Jzt6oJo4yQfrhVSdNNekNhQQxEF6YUh//EUwvJ
dkjdT/j/HLru6pmkDmynmzG3tV98w5hPoJXWpjXxn8kK1l5MBt5QBuIDr9lUXK667lniA8f+GJJd
73a9uy1uOBaRQqJwci0XjAFWw7vyRKaS/dv9wPgOEiK4PNxIPlFz34uW5K8W9paLnV8MhfNHAn1i
7D1El2UtmOvfPvgRURzec9jAq16tnDzgDQX6dnZqY6f0eiZOeIrx9xF0gLJratDWUvsLUfjMxX5C
AHASgNvBvuagcqbCAAQ7hBZrdqNuz441Oj4Hmjcpmk3Q4UsxH9KqXZKAftXY4VRD77ouo6SE8OHh
YRbxRSzBlN846lV+TkdAY9n/RMAW0APSWsjivsln97uRHQ66yfO+CJbSIHSzQCiNp1i5ph/IrUqJ
yvrDQvOraAReNbBVZfhSR2OALJ8aghcEYkF6QLJMRL3jITr65a8rqibiExLg3D6owK4Ly4GqG+1v
3F1diOG8T6eyasQ3LS3wRKLjiyuhC5xPmd9uHq1v47nw4o2dh8+dfNHmOTYNfNlGQRf3fcT485dq
FVoWdYM6YNTBFQnhjo6e1hQnqbttfurJoZ16ZQy6fR+syyhmPdfw9e4ARhZRg0HT0M34FPV0nAaW
WjPAKAH2ra4WO4338RMpet1snrRGRLUKawEFSO9b0/iN/qGeG+/H5JV/ZIOnMqjzfGj8RLfUZLu3
5Es+u7FF0is5AB/ySYTiC10lbzRpYcBl+iQu0KDU/A1JeN3FfBqczDGuTq6RDvzDzBrHRuJQ3sGX
6GXKpwaEVLSteq4spe8a5W5x7tGw9GWf7pQh3klCRCE2ycZ8dcUlX0L6NV0PZfgG8Qoppc1OGUo/
TPA75KuMRIqHWAJZKo89jvuB5I8FfbSN6yOXiSKsipmnMUV9S+V/cWwguCEYf5iYAsa3qaB8kVYZ
Bfw/9Pay1vf4G2oeQ1iyvN9qfPZ9uFY3CnUlNJzlkAFisMR+dF2l/cz2et0opUGeF9ZZdTT7Nhy6
OGH8xHq8AgX4wCBwLaSuzv4flxMwoDmKxl6mSPSmHOHItclGO2kg4miDNvACCz0vd85VNdXUqD3u
vfZ18yx7CZA2CVu1CKTBG6+U9ytZSTnjUO/IvcvUV5fD2OTvUkwymQ4PKKlm23WxSJOXGQsZnX/Z
OEX6L7JL7gapyLgLpi4SuCrm4DVxAUmJn/ha0AZNA8AspF4kjMBXQ7vX1g7Z8kjVk9Y6xCkr/jSl
/nctN0j3I+3Srq7YXSrDVpdKa8PUqBnsDVLEWyU6YqZDR9X9NvpdRMq5AL0kCa18BCEoDtZ+2cBO
Ku61gw331vwbylfYkCveXURtnIEah7Gj1VTJiIhmclSrPpOF6alTAxJEmGYPt8xIBlfNApscRS7H
RrLJ9DqsrpugE+M71IbvmR23od/9siN3th1zvFWAluNxMjQIMsDkCx9ZE3R0TybRjUgyo4DTJ+39
UEjTWMWLR1vQeV/ndJIPxTXbO9vKZwTPJaoXdV81L1LoZPYuhVgYiViXgtGQWm4iK1NJDAEK9/Z+
Y9s6pzfe8T5jBef1xgAc7nCOTKHsizQSIPB2ZfOB4zvwcHRB/6CiZ8jd1SKTup3cu7uTv5XpcHAW
oR469zjevrxU9X2rFNIqjPRwCDu1k1s6YLchIqTDtOvVAW8sN//83bJ1jM5EaYBRAk+e7Frj3eVd
ubvOpmrC2byYPAT9PJVGiD3C5Fc8bISc1qzh5QNiohkr2NkCtAEs/D4YrtGLuKbZPW2BRcRHN3rC
Jy9+foblTVv92sr38R2i3fju1dmRlzT5vmI5/Qevy/Y0ltI5Q872LG3au4feiIZc2r8ZgYnWfHvF
xMtLHAZ7G5S1Fd1Q3RD89ZcwavXHR73d78I0/We73a8ojJpfOZlXGQjpKTOYelzvlRQsIoOjKaqw
0tIm8+fGF68/wdROdDNlOjOjjlYA8ThFIH5oB2R16Gm9gTYwwQpS3JZf9ZKWR1DHavWDutXK+UXt
boOidZfHnvZJA1HXIAylaEthrAJj4oHG4rOks5koWK3dGfq+MTq4ZMkvXww0k/TX571CeVO1GKGY
mBg5VTvSVZs5GTuP2puWLPjUfgjsxabTr13O11IQ9sHTjS2YjxRnGIPVplmUuxmGZ4lBahDnDK6G
0j3Hw9h/+F66Rb28OMC2nIDJh1nprXABKX4ClLS1jCPVpekjRmxpJPmiNULIxNzuUKQnROKf376M
TIAwKDISz1lEZ8NqIenNWcpG36Zq1zcce/8ze7c1885FyuvIt6kdFagPnYpik6A5NRMiWcug4TIs
u8KPZ0vioATWaChuQrN1OeBbM/Pf69JfBoEqypUAm9XMRvboYvf78bUILAFHuHpXAEANwSc0wYOE
acQMKk88BGsIl1fmlFlPvsIiYWlrBeApfqZnxGx6rquNUWaXSs5FIwdE3ZLbFEHGeZhSC+UEBheQ
ZzDFMCGe7LMNR0CH83HuQnaZG63PrYpmtv1V/EfHyrpywbyG0NzVGoS9SNE5QNSe6u7T504TLD/C
cpPUcA7gC6QFa/iKPKY6/bQsSUb926IjG+VkumSEQV53XuAzMq2KF1o5hXDR2G+n975pZlUkxhzx
Nzz0NA6m0lZK/Mxsbe3VbxxCqsFmnPd91g9al0uE0nrIToJOqKRYJ8ia6N9LN5rExl8qw4ClMJbH
0ygcvFwG3nYuFn+BtoyAeoceBeNS3lYPN9q0sNxScfIEaeB9CjB5QDPQeml/KxBwRlti+GubGsjT
WxIys8Y5dza+C6tBFW3M8CnRBJn2yIQrcNMmg1Jbu1+Ic9FVsqFVVEOg9XKMrH4V5mvqmGL1+6da
lCEBaoo5lNJ/IvfyyAKNMFDNhO3g3C3zqm1Dd3HEeThAmeje4hqk+jJ2n7soLPon3B2VyWlBw94O
EjXb1ciMYkG0RPWyfZ/wgt2Tl0jsiuiFcFXgQaCCsRmUf9RNyuxjwu29WCAbefDbydSbhF2xNGzE
mv2g2RYFKkTQAfxllaWwRwMMI2wYV5K7xxI8ZI5kQbwgHemQQY4HS8NYubfvmvvyi6nVLNeoFPum
gzdQSO4qn6k+NQ1/N1htSa/6hq/bQyz5un3tEcysgtnJnbY+8fpErnWfeOyvkVYlykVqMuqBilek
des6arCvfDzR8DCOnihsenx1uqMYFYuZkorC2RAvGOg2Jjj8ES2tzIEBhynMBckYei2U9f3TD3xF
GeASyZD3ObgXQTcFqsFPb16HMfPl23uToqK3hrZ27GmcXN1APGpgUSOaaVYFrdVFXr/jKF55eFe4
22YQQM+BeqE48vIchkbXBXFMVe+RrcICMkUvX1HdzLpOrqSVdU81IUc4DTn+TzNaK2DoILAerHSO
Lw5wtMpOPIAD7JfhWi80TQavqugBH88QOBXskGXK7zBFvH/WsNlZI1oegltId6syK6YScbQ5CGby
nwvz2cL393fg1LsldFUfp4/mXa9mZASDkAqOBKYiI4qlLNX7W86L5K9WALcwhXPPtzSEFO4lKBSZ
91+ZMx4O6uMyDkUcPmJktLkkj/jymDgpKkymmCm+6cm/wpmrDUWJQBX47gZu8Tgm0xjCr3ZwGnff
e6U/0hCyD6I87+Ql8ScaXcThXDbx0LgYu2K/5Gs0R9ApSHBlb0Be2Dn94cV8AhDrgl3EjrTQqbBY
5laX2Aj/HYnkc7wm2Og6+sOjlmGXGPQkqP7oj7rxvHQsuMn1evg0gb60Onr7StheiQhioGBSD7na
5Z+2U9tnlp6NQrSlm2uAeeN4NgtaC74qeY+WYYacE8NpljnVhL5FkPZS2NWfuYE2hBAZIQXNsIAJ
4CRw4UDBgWDgmuUfyttRj+HKcCTdCykp0HofnRoXdjFhmWEHYn/L2k7l2mXEI5SxDygWgnQstIU3
YkyJ1VuK1PDZP+4K4D1SVbsguRV/nbW4AX8t8URVnWifsohTVVI7jPc1XmDYE2loGbb5vPp09m59
yq3NUo4Cu2yFY2jRrD6OIl38q2ZWA/vCtOFlw6pY0XrhxTrbwsfjKxUkarEnt0QcENxU5WdXE+0F
aQfhkEpQUjA3FPuiizpFNmWAJjmXNsnP02z/NKM86+Nm4cJyQfgYFdVKPz+sc9TUsArmXuuseFGO
jJNXBLmG9BhEzp+sMjLqOl/IcoHw7ROr5mRl7ivyMivhY7FA3I+n8cdKxJ2X+Mlbb5+pxSzyZVLo
Ko+Mvk9RphPSC9fIW2SGjQeyYWmAfy1UTgSPYBm3NP777aQhIDToNlAPQthCja8JQqKd7AGlOCt9
SSifFP4xLTKd2wT9A1mQLHTZIIv9MxgpdQPDSCAom3hXjdx5yI3QBikt7tZ1+wv7qVUzSW2OiMmM
1C+3Nyz82XZZWk187npuDnTp9Uf2dFTqLONXH0eVAsfz7/FlCcCfeJjKPML7nABw7+a1qlZflSYA
WqYh/E40dJmqB+fO2E9iP11ChWgJfxN8PQD+CRej7GlRdmkFDxQytCtfXTgrr4FcEwhk5x48VepG
jvUYiM8jBUK7T+00qcBaDDRBRk8wjDi+vOuH2jxjn/3qWDlygrl06tqroSIGWWWACH08QnDP4Ibg
bFkC+qo83SGclxcdknc+3xLSiwlzjI+mTncGq4iM3gOHpbCjP7YeFL0VFANazpRfozQsf0ilMvrq
40DQkm3w44+78E9ezUcS6Ox7z87xyWzDZIE99W6ZtWfVHlNX5OBhLxME8VzM3g3777ndhe5POpi0
uSKQQ9ClxISFBwCzbTue4x4umBa+/aDY5gHiaCrRYB3dsVTMV8m2WiN5F38vJ0AAdmvetfLk+OmH
WF36XPwLXheKoDWV5lc1V1lmLURawzDgtIGy5QUnRux/FuGsUF/gL1GnggXq8XjrD4Km8+qg5Gpy
FMQLET5ONQVwvUrn8Zw64IsEbcxfGAgVe9iLFP5MjrJySsXmBwzFbWC4m0SgHy7dgyX0WM2+yOkc
TzUfk+TA9wysRMFyzOKu9vZXbBEzmKQWtWqXI6nx4pPzw7e874CkXaob/gy29uutSITXH/sDcUIB
F0AU+/zcvojFPDzsj3Pk3FD/mUhCJw1EQqxkS1qId5Pn30yKekZjNF2MjySnwffOU6e5cJmjpohP
tLeUFh6r09hgi/mCYsnOk3RkjbdzzfE6XbNd8uR2QHPXOtOHDxJwDX7Yj9QkI+m6FE42TdLlpuRp
PRntU0fUut0g9al3cTUFS80g3KhU3RjJDqTJPnSY3fureTnbfDi3AUhq+7XvsizyxTldobfWFIIC
TBccQpC5uwwjp1MvyEYAp2oznCre4KjbYMhK/6+bBKDbWTNGlEokDtFs0aCMu/oACC+9slDOfGe8
xciHPgi3hjCLk8JPguFh6F1qbUZu2kE3fW0vXzhpeoXvsZSpxNZD3mxxUr2OASF03weKWVQ3lYOE
9WjbbDDANvAGTrnT1oPfNazUdXjG0owIgNgl0JtT0kEsivmXBSnUQ+0GsTvKN6od1FrvYRE5Tvsy
M7N5faUroyPeQeHX0J6eqP4oviTa0yxWi8ydF9HzpY0E/oyIUR4aK96p2hLRvUto8V4ynJXmS8vV
1Fq8Vq07SLIB55lw3sJfp5id8I11EZ/8tx/1izA71KoTJ6LeqGQF2ssfYWnCJbsDkRG/kE8FgMiX
g45oiz4hd77+Idsp662i5FEddu5v2cNuvKK3hCA0zaslbf0JTD4M79Z+/GKHVhwK17uG0UFLetVN
IWRIqkMDQPe1aZPgWaXOYMivHl/6Gql4FKBc/yRuEmKqe9/XBjC+YRTPwyWe01Lz5B0vOnG6/T8m
yQL3SmLzpca9j9IBX2RUTkYp66wjahyMLWIf5DKzOTiJhzstk8O1tSK1ApCsRX7zhPER7trkaHRY
e4M2+MOX1n0VulDs1mc3EtZpAoL3TjBsllCiYSEHuapTMkuab5gGbN2uCxJHk0gvxhu1YmXsHQXA
E49WSyEq3szUMj9+P/kxdjlNjV7d7Jsu8Kx6CAFT4K/a68wAQTEvbydIfqxxfliBJ/mz/aGc+21e
UAPpozMcch+cxgaEWHfucUijxailzCGxsbs+1UWaKICZNOoxYoNJWnp7MRWCHPh6s9Nb3YZsB47S
r5a0HulF1zrsY1TlU/bxkuDCCAiNXNrIYFQnPfwzpgnQHemMoA++ZxQWVbp+mJgMG6Jl7TsRYjBd
Vl6/B2jGUcCgFBpk5TcXJeTmKQM3YToW4o1dCmmrfHxvnfeo1z/mmwhLAVDEBr3l13KWLWkd5+mt
cckiNFBtBvwj97OQdPRIGK/57H4TWC/ObFRmhNS3yUzmra+WwrIsL7kAiqrh953GYIWVX96DmIGG
QufbIH1SMdKnc+VFrFl0uJ6vyumbnDbzwXzcx6swFDFKc2JKM0robYddPVrxjSQl9DGUNg1xG589
t5zM3QioWuDAVSBX1ElkgCCA76S2bK2mtdFt0rpk8pOlRxZ8b3Hol4Yb0N74ftYLEllE8xa8luTh
tB3E71Vhk43Eq2wHE1GdkTfHdx75Jrh30VroD5mS4FZqRlsDEpYAwof9QzvFLEPk0zRFUCM9DED1
BFBpF3PY8U5AID6ot0p1sOn/HKHTeNm2oBl69KfBqicFyjeKK8gWrPkX5RXJVZgWQb59dYx4uUdJ
8ObCu27TIeo0sr2uv9jmhascklpqGO7URZRLFkHR+sI6fDeJ9Pup2kuyzFse6NOJUJy/kV4YJhs9
4TiK0gI8UYWmqv0Y5KV2tquVUQ6y5bGSiY2XdtE/NWv8GZ5HBqXDiLl56Ivp9EKv2luiYagaVaih
49Qs0xFRNo+loCu8+Bv1jmk4liKmEqcAyGFF7QRoD/bpny/FAYICyoYc3u7F/ba5R7yM0uzwFjXQ
e6FRvSPARu2pgprDRxj5ZQlEYM/3OCMcQ68TMxX45q6jQkv9JpG8nohx07s03mYf3iOvknUqOcww
6n/0hL5weGjYe9VmtHmV9nCvLiI07LbfvH23HGNUbmjn2D46hqCC/ix6Xr/+O7nygvPQZG8WwTa9
6EPF6KhdH6sAejCDKhlvW4r5xb7jo1/fHeZ4MaMG0XMvboer7b1zMlG1nTj47rPACqAFLv1ym5TO
VcYCiCkGXSe35oSTQAKblKXeY4VkUlARwLIQlQ+RsKUGNpIBe8uZACx3mI8lKBFkMMjdX36Oaggu
SLetxcXWl1GHtzdnJgR3pd3NFcyEb7YuXAfnnt/n8ftTRaFBJl/yhb3rW+E0U5143AN4J9mmmWSb
ljVhgjfaX2rcuhe5v6my7sV6vjRRcBiDdT9wvMHrz9fTgux/tsD4RhQiAjR4LgPej/RNiiWdgkDJ
Zl+jkdkwf+icK1oHdjFigWi8JXP5ScWg9PKq1FxM2ic+3xJIw8EXb4KnRVpq0VYWdAaN/m8aZKwO
IyxgEvTNHYQDQS351yJdWo2stfMFa28eSl/fISNjiqFGuUfd+gk83I9wtDJV/hN7WDXvs67n0+MO
RGbUBBJb/8ZPCYllff5NOSNDl+txkbBCt6lwRvHU44QuECkE7x5zPT2ARm5wRqiqHjN3YrDTwnf5
pxtpTKNGm2nPoKVZ+BhCzBivPMcicBnuhZGZ/m77GHcnsBzMYaZ28V9y4xdrsRSGO2Zm/q8vuBFP
+GXeinFSWpCMf8x6+FJgenPx3HSgdQh9Y5b6to0u5pByL1ry6MbZR4xRy4kkZTMkxVa6PWH2m21d
I5CAasugaO99STNQ6Hc+AiJ2ni89r9dyQSS1orsw3Zk7gUNK7vxWm/QiAZhT9jPl1f1KukIskQHD
HD8y59VnYgll0Z9Db2XDEO5LBxmwckJGPdB1t4KNRbdOuqdniXFx+nmuDzygLovdhJpkazZnE7U/
qynQddOj4zdwhhyCKU+3epyZMq8FK0BXl9GB9ANtxu94MHL8kPNw6XgqvDW7LuNoavX7OmEVV8W/
1BB5rDjd3vyMnS6hphE3r3LkhI1qjprnz4IonAxTSVIoZCZ1ckqI22a+7iy+FYfNZBGg3HxA77Rb
byxDdUwAQc6UalR5zbMcAPznO1jTZqr2YpifppwXZEeMRWkpmH7LTOQaleEfbg1IEM0w/uA656ce
hpANwhiJf2B7q/QeUh3WLPPMcHONK9FU6MjBS8+m36wiPvo1Qkpx3VR3VXJDVrb2u/odvbXwP5PV
C318e/0loa3zWqFkcM8Oa2IDTe4morqwnu4b7NnCcit7Chje39XWLCd7NODFqpkZo3gY1Do367bL
J/L6zkDsxSZ8h/lh4x+glbUNuw74IuMc3zostkNAIeBTzzUysB/LWfw+Gvre8ATItgLa1tA5holn
NSPWh22RliI0xl86CdjFppfLio1wghg9mpalxdvCdafrdH8PoT8pt0CZtQV6aUwQYyNtnyfy11ct
bvZDEv23Xpp1GK+MHQb3yZSmCZUOQJRLu+GBYJeBDSpixdBICBkKcMVRZdEP4p+z842MlKEOXrV6
Pm+VoAbiy1fW/0EEa6IAir2P+Sx1Nb/FwYz0FAvrYCcM3WPEMs+AKX1vqN95QWfq2oPq4f2jsvie
DEbcjYZYQG93d71xQoMoBlJpk1lk0mzF8L0UngzXfEKzdiq83cPjKIHWr21QTiVL/Sqewk8FEMpY
U3cIYrsgYxbiKCtumSMTkFV0LAqyOuz/epwX3J7dUK/T4Xd4Fs4gv7aaZGNhlhroRN4tnJiU7OdT
GajBPY3pEO1Fr7HEkkD3jT7lMOApiipjqubC9ePHCLQ5wavMOTaQBSNKRTTiwpB+EgHHQsOS3YKG
YxS7udFzMp7apQmJ5WCtD6dO6IS547NKCfe19Oee9pwWWkulGz1PDVtRJ2pjxZlFKbfPorhxfReW
cE/RK9tMgufvz/PTH5F+MZbzdN4Jvq77bhlZuFdLqDTNFEVKoqSFTzOY4tTNcH3UAruFihtCOCYq
SwhTxY697FY0/+yYYZYWW1H7RtnMX4wQ7015JZ3ocxJGg4FA28O17BVj+RQfMnV6wUQn+GFAxATF
y+s5mztfRJ+pLgjb8TTmjytTfAliYuf8VCGBiZN8RrjStGSkRu6cORdLqImQntS7xBDcuFOxwyZv
rJr7O3FsEkm216Pt09i6VS9WmrXPY+WyCF3JQp+qcPehHEJ5rXh5FNW0yOse0Ltwl+H753KmSY1K
O54+P1g4hule3KMRYhJPFF7nRBKH6I2oCH1dEoFRbU85j8eJJlzzqyIHHdTR/JziuiPCx5o6gclI
hz3ODlUOSK9N3jqQyRz066F/pc8Vfr7cTicXO49Fl1Yoy3lmAJT7Xdmi/h5bHjiysK/AF7cU/Te9
1qMqg8hvYAoje2BTClYFsh2Z+Z0pX7uokhp6sTuOahe2IJfiK8Vk6H0bICVzPDGgJiPw7YWC+6TY
WVilAX10jbYiPNyv1bliXW7bwTkAVpn8jl2cyOhw92euH/Q714fSZ/lTKkBU36dynYUy3zn014Ms
rBj6WH2A32I8YL4l+Id6cCt7JP9geWQ4txJluiKL9Fdq7LdHyKXfyvtunLNQsPeDOQzS49N3mCIE
UNCDa9IrJCxcRRbIPe8+wQOmSDwkicgKxQPLbvrxqt/8KJl5t2FTM4brwXOdg4NmOKl4zs3hQPDF
jibGh0tKTgRLNYoLSzRVGOlQczEbQGW4/qT9YwjXxkswfHrvn4dZCzgS0bt3YLtUEsmLeTXN66Ew
3hVjQoc9WJwP1BvcOA48jPAf3zBAOItMUDNR9vDxQmGLFqDkRQa6hfIx/qT8hhwILvrGEjyfKRBH
Ovhc7kRmvW7VYBhsQ+SAdv3Prz8St9+iklsB1I0z1syR0R8VZgPBXIeVazxf5hSU7MvSukEQNhbI
Jc9nwAubC9WMofTCHpDXJILJyjdUnrfo0gHtHF1YBT7SAkqNhT+LHXWeyB9ogYcnKvIjDUymvK3W
qGWd3cHFjrKBgYvBqD1fgWczPjUXsCh3e/VETg9CfZCMOFTMyPDp+mMAG7CBO9/+qaFHxOXLEECF
g3OYFqhIU4oIsDD8Yk7FODdkLfA2XpTrcVc4KWs681YoHrOXbj0Lm3ZYsShs2QsUhheqf22yjEu6
kx1nmX++FKQpLuTfoEaNR0Ac/bZmZ76nP+I2Q/5nS5W3/sTQw7GDr7sDoOr4Y5zTx4reZ4KmWVd6
DxYMvB7apSjW8YkPHEIeVBw75U9xJkgdbxc6NcmhmGTNuOUznivsVAUHZsBFkzJL2jdsb9kW0Zf7
ccbgpQtbthbChwS23g8a2EtQ5L3moLuBVJSGPE5EcVZKvWwL90d8Q/CFNLojqeUXA0c+eGEyBy/1
+0wql1KL8iek+aYQdYAYa8+iA0E1SdAuYCaIW3o/HA+h9sBPTngaLR2Yn7/Xjbe8KsQGYbIrieaJ
dIL2QfVzS86POATrH8Br3SqLEClM1x9iaUggN6MPSU5nDPS/kMtVGXgst7d//Az1ec5UB8vmYJHn
J7CIyk2juxC4vP3DSqGlwONCaSO34qx6lPvkLzGfevh4tqqIiVS94OiKP+weDXGsjz+XLVQtPMXW
0v9o9T3v9BWdYgHEZU/QTTv50ga1NdzRZBd4gsZkN/2lfwFCjpmEpql7421rRxp4Gyd0pm/iW4UW
YhlwzyEwBdiE7p/8FDniTjI1MOGkHwucvsVT4A91VHfgm+wzxSp3jmxBojxYt/vrMUxg5pjL7IZ1
QJ4jkiNDJgW/7uES6Tj0tqkqf+hIWXSxeQE5M4hqStc00HfohLGksXh51jvVduL1HYdJjZw3xdeI
xhVic3FUEAS3jvgZMwK3OkDL+HDoXDr58P89W1bsBoQ6t7zq/9+38s8UdJHGTAbq0mVdObWfPitL
UYjhmxjXU9rVZVwLYGht2PTmYz7IbS4y6jHr+Tj/fO93ypd0FCGB9PCLsFzcUEFI6ScaNBt63H+V
ADnunCByEs/XhMpWoV41WDsZiAXbOC7ripiXYPVgcdI8d4OYJctLnRKrQ4ZFVMJRZYtFOttekmcS
DdrEeZcbvitftHU7x/F5ENlwitGEDblFpzaqaSq/4XktZup4kC/pRB7HXqp2Lfz0e4vF23foX/mc
JsnvgkirlJUbw0WsZErflbwDBx7sSHvkLEW2MQYLA4op8j2cEgWNky9hdXbvwbCgfOVtMKV/3bCn
z8uHmnesyO98XULNSt75Orm/DGiy2jABYBdc8K/jYdP/ReNDZu0/vy87V2F2Wxhup5X7iBDCXUBI
03SWootH/I3rdvx1QI6tED7XxPVOwEr65uhI+f142g3bleZQD5+QfVBxl/pdTdx7Xy4WsUugEL6W
kNdfMfFdG1rhnIgiNmtUCZG8IgiJCXHu2YAFFBIgHu2SzX2/UYKkdT10+NpNTGRAOA9E15T+bDPM
dL+w3KkIk9GG0xIkC/qGdtIK8/SI95nef9VvMeSlNUlyqdgd+wfsv0XrD+VPrglSnDfMtMFMWzXH
iRqL1/i4Whx7Ta8+85izOLgJvWJbDp9mgSPuTCAAJQnc0G29j5lHDsbIPXVhS0kZaR1uWM5xiWct
rAtL43JlTadkQUHrImiam6AdLpT6v8R1ud/cG1Bzh1O5RQNqFPeKTXacGzsyPnCLaRzHnm2aHJWF
hETY+rLAAUhSjbnor4bk6TO8QCGVUZ4p7xB7XBwlxwdL2ZXwa6yD/B0g1hx+vX32UDkIE6PNUR7A
EsUsXBTyBvsv+WdwCAugPNm65ha5yJCrvUMNWEf3Z7KH5F0M/dI2aP9b/MaeA0lI6eWF2O6aQvlE
L0rBVtk90EuAH4IkkBSJPOvC7zoQOyox9aregpZRFmS94QORfSbW1vacqCI8kNpWaqCylx5gGvkO
WAghdnFgfaxIxi6jsTFgEYEZYnfPzp+VTmXWP1K3sNqjhU+iNqXsSJYK70Hrjr935/qmbZuf4ciA
DjnMiaLNQCN6tw0GqS9kgqJ7yuTbg5e8k05WBje2EC88qY+LdeWFEXwjmJKrjFkNE+Y9owIxtmFl
i992eegXFVrf2P+mJiEQJeyhnChmg72xV4azfnAeXVUqvijNtIM8YjLOpurMaRp7/HprYfNy/MKt
gnfyhd+03B1t0gzfpca1pjr3WqfSWHfB0+IgqTVlII7BZqssM+lU9fEqZhKk7y2yRKnQ9Oi8eUhr
0te8ds2/UQudva6hb0mreb8m3QT4ZDIFVWjCrU3vWDqhc7c0DDHxznrSRo6H2uTBOaNuI2Hla8l1
LlK8h0+ZMAPwb16QhhP4MSPPYlLuQ0mKg0sXGznUJciq4Gi60EOGAyM1XHho9D/kc6PA/AJcFV61
NCtrTqpLzYOzbNW7q5LGA+NZ8wBSOsmEWpV1k3S1Cz2Mnb2U9AfxLA54sXVlzfpixMKGJv4CciKe
NJOmYyoHNr3Fp8TG23uetkKSEZa7g6dXR51SrBpn3Qu4ELoxSLE4zP5RnrYIwMA6aNYaDrMK5Axp
NvxCGmEMFh5QEelPhBJJrrCOu3tbFe6XzoHXeR2ITQu8rGM+gY/p/tnm/MOlcL76X835U8a8JOdB
0WAJwl7lNMHpFSgHd+pScgCd1C7637mcwyi46q9Mpnu+9/FQZ3J6785VXbQmuyeeePu3hlwVw0gt
aqrKr+w9xFnIV7L73eHmG0H3L8MRhVVttL5uq6EBscr+fVRDmd+XuLNzCMpFLlI0Y5woMKAwZK16
Xe826F6Lz8QhF3/ctmcXzI6cMZ8cBiscQgq1koAU+UVauBP/R2bSvciSTH43HM20zkAdXa8sSVfC
5hYB34plAXDoN5RFnORX2KSC5yrOjBYlWkYEvJY60+CskEyLBct7hQn9p8UsfeTpM7LOzY641dc4
+XnGH1KnUS9Y+ohJefH/qDmLLtb0kV4OuW7/RGBWQQVDEpkvSSoCahqkp7cC1TQWpHSK6TACYS+v
RiCgNsmuMfTi5GAsJ7hx8DPenkz0+Is7AoDF/0tuPz+N8rGlUlx4c7alXCUsEvP4WaIwtPBeQP4r
At/OAs0ekUvQL0PMMrConO2ActkzsBD+m+F0hNfaGacp9jiILtEQ+ZTMoNM0RQrkD5B5ovOA9cEX
6zsDvfOXpgEEuUCmAOO6chwYoxEWZlEOG+BVzTT4pMMAJEqgaxyBy6ND5DTQusY0c3guxeUXWAon
UGVsH/7jQLzHpeRzX1SJFfkqTS1utPeFHSJqgtOtUKidWwHoucvCiS4D7uTCc4X5xsLRJGuh2Lph
2j3Cs78MqFDbWNv9q8Kym756sobdDXnHZuIkDGenN6cdD1jikNAoMeMG584JG3HXrmSxTIJ6D/cT
rIcyaOKhaBPDcNkZQjJbvO1RIpGvq18dndFCakaapMKbkqeejMyZcpuWZtW8/C7esFwaM9G/92Mf
zq2rm0vlA9LbihzM/1FHguHgQIMIASG3WyO0QhyKlt2ndeqro5nD3VfisbyGPT1aqRnrhuxONRYF
ag4u7xGT5q5Ppey1LTzoekdI1x1lXesFyuSkJQBNjgHSwOFSK45HlOzVNcA4+EJuUnuDmu1tBthR
FjM7QPUNBxB+UiW+CNEZkjy4paGupV0tIU7uN73Ki/B4O1eHHAmzMqWfXAUsHARgEkRiL7XQQuxa
X3W/xQpE7OjcssR7jFAYgQ5XC+10DHXLHTal/4vLBtqaWZHxRRKHgZP+OfwoMkRQjnwGwtm3sjF7
1FSvrplXJepDHTyhNkg6diw8jyuhtYkZfkmju0DF1yXhnZoPNXn/NWfhmRLdaScxVkGF+W9Mc80c
VpecJuStGG4BLOcDmOnWcR+9hLXP9VxddyQn5NqN0JKge0kfPVUv5uvSqP6mN4C4OYLAdzOo6Bzp
qA6bG3hldCGSvZf7aVhFSdWCLVIg3FWOPZo57t0GQ+hbwInQBP/XC6OHxjZgYtbfHi1tR/bHgYZe
y9Kysk0aP1j++oPZF+JmIELecyXwH3r/2ampfnvGCPkQTAlGt5emKUZOXYsgms1Rtuf2tiedT2Fn
vLaiuOvBuH2s7ZWczgdgc5yiMlpfRVTtC9KtG/s2K0zFipb8Z+e64+nvsCA2cmfr3IfM5VI27TJX
H5cErXGNygNQQx251M0C+1CzCFD068zJHkdJyu/OWCk8+u720YcGfZEWtdFA4O87E+dmbdDKpbfJ
YlJtvoNekb+oIttiZ+gxHw1fb+EnkX0+/X9L/52MHH8AdfgV0owtQswnFDCwYijlqiexVBxcZA6y
0k1IBUqyMDYFn4TScooJKHW74/JPWNqZJnUMRGKZZZoAI+ZXYOpW1lsH8QHO7YD3mfEm4ZFDtMV9
28vIGbmtkF4wUjW7+q/TL5gpjC225Rl+nhfWnw7rHJy3V28cPv9zTgvOWmawJj4PjGfFRqmBMc9D
ZbpEmiDMP90Py68ZKqWdJ0XTBfVg+tN/sn35V65YS7YogkRI9sCB4wtSIhni/L5zVcFdr858kpUS
Vz7jpysGA+tJuswcriomQxOnrgSzESYUYtgKhx85gc7CWlXkAEUnzBKCtcQefviC+FrEibPgMnvw
Js8GvonXmVt/uRDQELUGcdgsq1bBCyVpOojOBpoS9eQGbEI0oSaaVbkw+BG4dHdPZ/XSXCth/vw8
SC4i6sfRfj+Xa8lTNZpEv8bO1YubIAJV2jZaZlOMsyaspXVHZ8wZNkjfMLdXqAKQf7ebCWFM9/eP
cJteSLOHvfsGEpbMa1M1SKupaTmiP+1gtF0L29msFSgrRFoV8CyxW7uK4u+c7vHfgkzC4euGOv7Q
8hFhaC9xmtoKtVPjU4PgLSLWV739Rln0+A07RQ8kQPMTeGA0yScwAAN7xHEfIjl3kSPBjwStcGco
8IahspMCKRTGP4Ex5aUUOsz8Vih95y2Wx2dNMwfuBGX+BekoJgfAmZeUcg/X8ffkUCbGtXnmK81D
EyvCXDOE8/O0YnauDgvQA5vPGWHCKqOYV/YAQ4HL1GTNUGWoF+cffYxaOPZuY2zbEg9fGfVTkMd1
F3SA2ZORGSfxseVyyJw+CNl4NAq+LxbA/uZnMZ6Wvk7iCd741lx2ek8eZhL8H5yAPU6yftmTb5a0
8oBtwVFm9Qb02X2dcXZu8M3YKGmr4a5fabvB0TNfyM9DVMrvQ3IqsvlmNbUeHbJdd8fRcLucg51A
M/+ZNxpTmAqPC04oPK2tImyPQpeHw6dmYN2llI9D0umg24vO+oQXjGeh+0VT7P2VVF1xz2cfi4UT
byTxRVKdljRBn26lg2PE5qD9+Tg9Sjldg4yiExs3lr1YL8Jj8OcUkAsh780HU9VZddW1CuE6fj7l
N1hefCNuMeBpHpuDFkckG1BS/UY8NYsr1q1f9AF9fK8kMbMa63mk1H2+8C5SD9YfopbG0Tm7vTh5
qQ1niaVWDn7w+/QAP4fEg9NCk/cLqTx3KV+8V/6yzPDNv3e7P8ZzWIZLQD+AVoFsPPynvFa5waAa
WmSRXgHENOnx4Xdy39DHMjD0Xz20cxI6TBf9ejAZrbUQlMEFiluDhaOxZIwJqTcK2O9nYx8Kvz6G
hkmA9c7DroeAPnZbANqCtz/k8pfz78ml6bC/GgK1kg6yUskRWt1A0re29KXP9F9UbqUyQ38xPKfP
rrzeIipJpCOzOvJjvm5h4+fzf3irAoLIYc9EQV6aD3KWtcatnIFwtMJZ1XqtTkZqj9Bt5GwwbxTu
4gDngahi1WPta0/tspuxeEEtrAmfCXr8YN8RQ+JT2jyB4/sRnXEYImOuzwQtilUwK6m6qNIbGBBr
RHZx+e5EUx30587bI3q7EyvXoIBhJJXfy1de54YaFlyii+tIvOK8skQfGU0pZ7jLO7pbPTT+k3Tw
VJBdNxm0ZB4a4UQY0KBkVCo12DbKto5eIwnKsfJnEyp6IOXQqo34U3UkVZDlLLTYLMWwQFHiA3Yf
tt4z4EynbOR1zPMSBVaPmnyIIpVbpgpQglMTeE0V+3Nbj4BZsWlTQ4NXTBQYq5fQGBUid1VT3cHC
vE9sPYtmqhsr/hyd6oFbUmk7fu/H19JtH9+7tduh/jqPFvw2GCzK/UmKJoujk2ZC3F1Tm5iphBzS
Sh27BTUnE5qdqJhDMf+eo+3ZntJN5RBxPlkGz3HDWOGD6VCuzGU/nwG0FG7KMNIruQR3Hjo6A6+T
rOGjxHinCD/OaBgHMaEXragsee28Jx7z3+lXkvMHt4VKPw7okxcCbzmNXPyFjmOii5iwYODXTypG
J/Jber2bfW+s+Ocl4tM+MC1Dq1FK2E0HMNAKF490wnGhstirqRbQ+iSg1/Cp8QsH+IfMM+b2B5jb
3XzwQ/oQih0hNmv54mNMl/Lduz41tEO5XSUisVvDJD7b+KjaLtzgOYtalTsMJdgEgXSmhLzcqR4V
W212b2bFKM/ciTAmuqbkiTbB72nicRRdHRLpD231m777btliJUt5xw3CxANLfQ03b9JAipq0Yf94
+5HWoaXuXGuz9tNjP1BgbjIqX/YnqzwnQreYeb/OLAX0bkDh8VJU/xy+ZrA6AHB9sQk3t29O4z/7
qBkfm6DgxW6RpjKk3Ua9zkasxScjXZYVVkJtnCMrUB6MZP4cC9ABwzsRxHz9ixD7wxM4LG7uZ0R9
lx4rY/Wj9d7ImxLZReizFuWxMlcQlrk7RV1fNu1c6DgfPWg3dVjZgrg57KWDMPLLUClTAc3Qugan
SQq/HipW6OjEZlDuZMMj51mjQkUJq4hgXQZ8bJAOJrPBGkAfctrPg3LN5IMQW2OjAtcJzx50p9u3
Lfs5VuPVdUQSJNh4Xct06T79TnjN+ZsaEMdrb1/U0T6wJzbOrGXISHcSlONaB+HIeki4tuy7oc9Q
Ul6x983FX1yVxRFAjyWiaoyeq4SMzfOniOPSfp4VZvagpdV/vyYG2YmvQawPppPz0yTo+IHChWOF
OEb3x4qXz24QCyQaEVjOSUkfUpnJMhYorwIo70Ewq20DfYNDmBzQsBDnMRTuCQE7PAOYpxbRLGWX
VxYf4ZLQp4HZ+VlF6xaGgr4bh0MshTjdsKl7UnnVszxceuNuZxsBl9JQCe5UyY8tyQ06FSdf2PF1
fD7d0Z+Dp75w5sx3TbeK0QLfcA5AtBpc3ykknvwOAWe7UKFZrFRRIBMgTa0nqbxNkoloUWW0do9G
5Rlp3o8Y+2r/MHtP6eHm/rD7rslVfWPtglEUtYe4Xn8abyYx4AAq4WuzPSJ58LDN36AKSIvngZdx
bl8sPbMalDwCnL72H9/2//cm9FL4Qo13916bwKAMqaN88XbKSsvRFa99kwWvteKTS8NwFi9PYMMb
Jgjc+tD0MuHq8p415gjD5VQ2hW2SKEwE32fPpcQnD5w18tYgbN+8ylQIYMwOzjFxzKtZGVxr2jPX
X9344TUZfploKcdJ/NDb7QPjRLEKacWRHfHiRpx0K+H6cFr1oNcK7Ah6oMYgLRwE4us9APXS3y2d
IaA3vQ6AlWtqA5CnCb9NgGCglha3P+XQ5wmrC8dzx7Zh8dL7WkGOt/gpG77r4np695ddlQOzn5FK
UZQHFVZmhcfXATsHKKcVHPqc59GqiZasAWkanr87TPP9OCGjWv3g9mmfPI57mWMwmCsF3Ja9Kd0s
p2fgMalqzhvccHO9zI9SM+dLd78FSZr0lMsYWDxRThAuUSiWUNwpPiY1wyNDOSq8W3PWAW/X/9mZ
0nJC1xWTxqkJGTgoF9KE1NNJO3DO3IwFF7jYS1wpMItGwD4HXpusAFCTuU/BNUk5cqOID5dvc138
Cm9ITmZITc6PgLKiUPCFJs8pwU89Z1+GLmv5FLpJ15TMacJ1xkvtfed/mhIAP09Gke4KwIuaErPT
dbSjO4aV0aiWqWK5mWQsuy4pJ6r3W8kko1KFCg52k3vr0OUDsn5DVt5r/dDeVAUbzNbHxWeHPBoq
3j/qJ3w+7/0Wi5w3N03D4AqyTE31Qg+PHdC78ydb+eXly//2WpYV7tBqOiUOqwr3XMiAMxECuvtq
rIhSiCMZ7c9PHFtxIewCM+JGQ8CC8kg8rnfPPjoOwae4kSzWxlCyd3GeD6nlM8cBBuKdC7UQjRTZ
rdZZD5H+EF0dYCi9LEt2fIW5m7F1siHeA582ZpBXiNiC0rujpd2qNMoKgJOssZ6pOVEfKlXi8qAV
KH+dr0vh2URBuwTGWILp+YnGxe5dLm/EKlxFOJBhJMgDBoLbNac98bZ0VmXFRM2YKWur7z2VSoZ0
Y7zQl0EQxLChs5MFxwDBwju+kE9RDRW4iHK5lL7huhOretIQafLhKJ00eVftrOiztotEX8UHs1ns
DLuVgby8XaO/xl0o9aUmiC9XxcPoRgLSCWFv60Nz3rgFQ8f2NGMja8F2kfmHlazQttP1Vv0LhDJM
vbDSLCOf3+CimRZX5xyuPoojtcQv+5DrjQkZGTRd6u4qelpwFlBSI3n/N23iCXm6fdb4Di9yMvXZ
Wv3PwxHI9j7Wnmmb0WZy7WRR4C4B/QC6aojqtYszL6u3SZiy+4b56wosMeal8dSyXnlwv3wYIfcl
U+spIs9+njoc1QbH/7KiI6Z1lYmnirkwzYBz1aKAw6IvnWSwRBB0gdpEI2/snA5nrpfmEQ2xH92a
KKwWrbPpVGGu6w9ma7WcqKtkZ/Xa8QoBJiJP7bEJ5puiy/sP3d1tETSjKzNqTaQdVo0dJmEAF2zA
lolNNXfPNlsOk/Ecfx56UFFCsAW9n/EZaodE2aYxGntyd5TyqUzc46KWzXhdYQ9JkJ54O6QCF8K8
W7wzKDEiydSLsSIFnGqjXQgbmeV/5VSfuTjHd6MYbRNLvoN2G22qXOp1aF7Ch7lVF7RoW5PKhIWl
cWR84TO+gNo0VcIqY0LQL2avM444eOdrL5ST7BWZyQZ2AMmfX2011sZt9SAc2imy5hUtz66a2AmW
aolCEguYV7cDupbt6ZAS5ytct/ndYv8YE7t5wl0TGojwQBbuJK1jUPXC3DI6QWs8QBA6W3190A7c
M/9FCPnZC18l6TWduv0M2T3jAwLMe0GcWduGQlflZ23lRSGO+/47vZQga6TzWskuC3oj2Jg/DEHB
kRf1/JqBhACTYXYglsPsWyS3uXA3CAr8xcTobABwRuLZomaejPscgpx5/nvENsFukGR+lbZHWBMY
HjtWkLeh6ljZk49InyA+WU/2cPxbLPcSMFKJfN912dNthsXYT1eakbEYrtHarZPQRKt9bi+m77hk
yTjKd4KC95amQ7do5fA+MTvT7vab0ofR3v5v22rM0+N6hX55/gjzX5KI+i7xvMbeBs9OgTE9rGNc
kxqgUZ7YR7bc4Bi+DTHVWLEH/VWzCGwYJr6+H7Lid0tnZKVG4kFRxMFrnj8SC2OiX/tcKf2PqyGe
Gt4EZ+Cz7vqV5Ljth2ReW91HpJBFjBF3FH8t7mzan+8RVLuedTPhs9zCFD2JBo4LuwwAzC2n4WQF
n1cARr0WG2yOfiAujcGYUhHlHakFR0VTJDT6YQjmUxNgjKYAjXZxsgyOLJecylcwBNi92sx4LwJm
025qMxPe8MYPjHlT3hHXDEp3wWP39f9Y0E+cP2ZsQS8LQxuMd2FzjVoEkA9vPmiGsxk28DZCnvaZ
Cyc4dPNbTUW3CGJqQaiIDt7kO0XWAlLy0aTIVSKklK1l9eS56qa+sU/KQuVTDgXdG+rB/pdopyxp
nhlibjyntLHj0S968rca2YTZFpfT0q9kZ+UykH9Efe8a3DtI9W4inNnxpDW8HyYnw0N5eFMJImHR
X/0S+nSDvHz1i+/nQEju8PlPvAj2xLKbyCibmkwoGWnaSLvFDKQXn8SiKEgFeG174hnchQsHTOva
efRJ2lhSH9QlmDMk2mtUx1aAHMGsQFOk5WKox6v/j9y37huMDe9KpkiE1wFB/hdyBmcs4wUnGrDE
7P9UYpvDw0H9u2k6rgNUi83FtkHqAh6aySMBLyTCN/ea5g+KW1G91Tks95G+to2jRmxilew4Q1AM
rXVAeA/++0pBfsYUOLEKraDSBu7pcy6NXaM5dcUz6vnG9kmxmmyi5r/qTdwkBEUp5Lv/LiRKfKlM
mKI3CAk9hppr8ZGPyX5ewun4MbxD4EztmRci7QchXV+ZIE4yJUUr5903W4CZhH0562TLQhyHbK5s
/KAx3JYCQchhGi27sqIjuBk3uDfrrycbb4adlTsMY9gt3Q0sDgtPu0Xlu5FEyELjz7lFoygYVbUx
/2OHoZumyxDIb0JFaikynlQwl7K9K8GyV1Qvj7pVKOTvNKHjkH6OTf6Uz7fpsgrME/9AAeR/xAAi
kCYOUKseiakSVJrR0Ixlld1a8dOAxzlPSxu2UOYjT10ajg/uCFGX4dsFuYSOQYopCHPkqgClPg1u
3M+jNJMgSz6hiNIrfqqV9dYmSMTxplfC7RGGI1OPqNRkgrM0unBtaILb5JZ7sKLEhdFtYeHFqDm5
2T6pHvl7HFIh+xnGhQFGbHtaluvl5av8c1lj/jtLhkvSMmy8seEY9RrfT+LzErHcFr+3tBaS3MNr
P/xLSMIo9BB7HtEe3/gY15xRTl5Qp47CyC8v5gsNfoqQIRfCUT9GCO2MOcnpFEP51uH7NR35sCAJ
UAjg/fk7j4Hwl0H1I8a4WgtK+dcsEYVbpYdzu3qOvkgJdIcVKRjp+NrVbuoklCULPFBdaUbPk8Sl
pRpvwS4boludSBDjXVLeOssFpz+Np8kw1dqE1f/9oVXOXvg1JC7HYTmqIzXLBkF3X6WGgXJ28Z6s
NmN7jErSVqzwU1WPth6sHbX/oM2/iLCGWCeEqOa8cDKAmG73hQT2bmNcK0/PUpPHCvP+0jpsoJ6w
M6bev6roa9YDpxlr5XZHW+SSqi4h8ufS+rk7gtXN7DBPex23scO+nk3+O5kxGHSswZGvYgxktzig
7TsicsCaKdVlgeXT0AgvgfBJB0humYCC/Sgvup/sfmvt56F6V/1RAJMZhwMwKtgHVIiUVTbutrVH
YAVL56Hc31yDxhRBjDqyurYG0TSI7b5qrGh+SnAt+5B9xEnTGJB9n+DGW0XE0YuREv/GO+Q+XJ9z
8KBaqA85WTXf1KknuAw9Pqbk0gN4SjLCEzNnDVEHQOhaKg/5JCdP8hx5bLXm6uOBabJAyG1BGSCG
Og6TOEDSQ+viYcjGx/YAJzY8nIHgCnQudLdYtIa9C4I8MC+rZ5RnQ+yinBVTXRrDu0y2Oopxl6LP
YbtBC4VuVoaWGhaV20GpZYCj+3jTqg9vOCe7QVoOebyYJRIUL89zrIGmbCjAUygD0XBNrdQSEwwH
Cqw7/3HI7wsdUpar9i7hxrFignpbYOkTF/HR5wSBW1dr7tpdSN0KC4/3gWUvRV8bKvRxCh2ICcHG
zLjHU2YStRTpj9iFdpg1CXeQUtdiFhPa0sc1HnwtqNyp+1VSIhoWfKvc8se8xA4yxETXISEKV6QT
Qem17f4FvAfUI7W/2CHkaf9Ua8ycC0Frsb7kMy73nOWUiiMor2TkXCIBy6GCT6WfFmDHFJcChCaK
hHFyBbsID5bKC+Ga/qcbIt/IxOEZ3maVckQNuf8EMVI4xB15Qw5hkdvwIOGBYzUpkjknTKcKkYj1
bXYoV1TUR5i2/839NxCUrCyMKM6gAeQS72NWNdgEvLncO7B0IYtOrugbeGsyW7DCbN4A2WEQoRrO
Yzn8vXOtPUky4dpdovd97eU7iwogTVeII/rhEe4LPBo5j28z7NLG7bse/maEl2u5sA5tjrjuCqe3
kroxM4TWmRaNNL+bS97my5oS//KGWo5bT51S1M3pDBuQ8fv8ZONL6thx2nz0IHhFt2Su6tAfgY7/
alfn0GVAKxkRli1aplBZ43dKCUGZ074ha0aw3nynKloEFpaZSwILGNHLzQosKO5bVn0lE0j6lhLg
zUl0Cy/ybt5E03ICmuyG4fE7Z3cGBOiNZYKhp72ulmNvRxC0GGXL+C86cI9g3JSBy2aJQPxQYKSC
Uzr5byIZHpmbs2NW+yQN/bRW6sbHFdJyoX50KknjKSYumjbNzi0fnDTRGpkndr/i2BJPJbvADXR8
C+gXIx+SfRYd+a1lR6ZLfl4OA7fgYYmNkNbJ+1ne0K/LNGRmNLFIDCp7fhGg0PZlEb4P6s/+ULwW
pY8NHQt+wEWaYhFtGNck1cDC01ACEXA352wXmvSar4ZQ1nFOLCUxgh8kQ8dnFHP+ffWdh5AXduUL
SfvcMOKRsxDmMMoP4H8qIraw4au+GB2uGBVixv3bocLA4tCzItIHDmhJcdq90Nz7x3rMcDdQZblV
9VAza3Esx1DK/X1JjFWCjiJV0rVQDBHQkeQt5CSmcG9nSSBfITQjYeyV6QFZpStEjzdjPqJwgOej
dGNQihwZk0mE5GZTZvwK7JnbaoN6ysFihxCrJvWzjPvcLdsq18/+dMBlpaUNmcq695//L0Hcke4m
J2eWn8p9QmxTVU7sGi9qbnq8gBSJF2AlIeHmQ62oCwKTySYVnXnWtBQ+h55MrgpmZOS6hERGUHuM
Zgv6XV7F4vOkREiDYgMRQdEn4MH/ucC1eLfcxqkD140Ysc/h140n6dn4vZMA9ZXgQibO1J0azTM9
VWFzNZPa7xNS8CXUjwBTXeUWsgjhVf3DMaNESUlNUfLWrPzsxlZTnTJaPMcYPgvYok9D61Ao0Uet
JMY+IeerSdMe99ciEoWEz2sR+MzRGhJ53xeFiHW83vPJsheCqCr9h63yco2f42xaDMtWaJWeRQEs
nj2YHlCYYrwIbu1G3xMuF+zY/tNuDq/fhrPpCSMzcmKep3sie8UvzARAJQalqLGP2e3lBzSrFc5U
dPIx/yo3kPPkMtLSeCRfArGPYNo+FM/kylTeJnxxnCmcxWhuylUbM2jhEvbmQ+hlV/oPNsb815pg
zYL5cO/ADDt9XqPT7z0PT1Ie86XUQmD0gTj3BWDh1AXgdD7PoaSZjpWzp93ZABhZs16l5l/Lb+zR
8APDPhS53YHKRwmhoxjcDnmCVphZOo0v87pdxnHA/uP3SW5aWSB6GJJ8v+5HQrlsI+fDuZsymQOo
vlhQQYbzDcLYhDuaIrCJI0608WJ3hc+QvUs3wtUvOfMjQTUdP6yc7WPGPe9BnZo8Rg/twvbCQFSz
1Tsil47v02c4V6756S7kK1hDV9TASxsPr7vHEQLLwCdnP8AkBqLvD0szxfltMQLAFVJv6aiHnuq6
XDn1H/5jAZZofxxr8XZ4YT/BaOZBQJE+mbWTphNTUyDMgCLgS7SNcItFmdpddYG8s783eJbyyoTt
zpN+aUzdabO/Tm2D0TSRNbKLhtWsLyMSRnr1KeciUOBpZeK6iamdiOwFN57S0tteiuMLM7712G1a
N/yCIIBHk5aF39XyxFNdpV9jJ0fz9spfkSdg7UkXqJpD017Y/A8lBx1Tm6SjwnJ3lQp1Z+e3imcH
s/LOCwv9KvyaAMaIOb9s3chzvaf5S85EW8VW3tW307flvaXqA6qtXxSPbXtc/UTscyOY5ltOVLVE
AvpUVWMnZPHKULSJ0ppHeH7NDFpGVR8GoSvXfbMd+N9gIhLXAyoVa7JP+VBokK19mreO1OlyX59i
yW+mWRGhCMLhG0bapD0xkaBy8PCl+t9b2oMzZd4Q0Ed+aWZe66oH58VETEBealiL24V+BAQpNlJr
Bia1No04dI6nJ9b0pcZHBxrWEsNVa3u47wrfev4zJxAZ9Mc7ayo2bjXzRs9DO48dnbXLNu58QVdl
lDziPD76z0LfHBuvDOia2oIfb2FI2ly9ebMtRsg031ERtq/9hhVKsj1SsBCB532BzW4U1OsuwTUa
j4ZChBgVrI6mxKMAsYXsLzdjEvFa3vWT1BE7Z8s4W7vYlcJi9lSueA1RucDlb5m9PgJRITdkhIWv
D4kXIvNRrLCVzL6u0R+gT1M+SR1cCjzvG0QzqWegBYOPsQMU+y6YykPlAG0U/aO1Kglw1TY5igR4
3VsLoDMyn9eJaTzPqk/J3MQeONZe1bZHaubqyFVS90JtggP8G63No3bqoWNmLbXubGr2igwoz0hI
sD98ZOlz69w3BkzwJomQ+LaWGp+MsRkOcmLvOyWGyy95vA8O9MywgTsuOKrSFeztK27QhBz0/G7d
3MVZnzBxPfyMklIghI7k4//tmtFp8ECdb8xnpgOj0duQSfLS1UAilnMhsGDgBCYFv7whVX8+X8lQ
u9dQtCnqv6jhFLaZnAYjgZgsSTpThFDzwiubaooMXX2+9uDzIB/hXs87RKjoze0kM9TmGDYMZUGv
psQLpFx1ZOrb/9ocjx2cJcdkIoZr/zw/ua6iA7JXITBoYr8gGVN6G74L1/IKGGznOjmwlA1VcSCH
bfrZiKf04JXmb7VFKVS4YyCj7PEPQsxVNgS1TK910Ad2XFmrHNYdpyYD2FsGKlVVeoltoTQYdpuG
C8raybnoumwdpE+eUh1ZTTacQHfZwY/qqhYabmLSv2FB3ZSqVUaj0hSMdcT5ScHIvmpp0Gg3WfiJ
kW9FYOO5mr2DNLnkTBpKckfbGnSgKYN27ZzPRL/0dK59j6gaRx6LS+IqCCtKwkhCPoF+9CKH5z74
4hMOCgzqk3qZCX1KKhP0Dp6sBAOpzdf5Vvtu8VrjzYatWuotKPyEXAJ6z4E5BjTfJmJRmgIF20CH
65P0zB032CaQY676oYZGV8jrxhfp0VEBIfByhEmEwte76l22RnVvyPEcClPmUI3QXW0H1qmeU4XD
6FQ5/hnPR8w9kH2ug8TL+NRTa/S6FJhIkTK1cKhC4yCc+VZ73qYqPlpsu2r7E/1Bt4deli0RxHUm
e5lUjeLFrgMCdLPf8i3XQhWMq1mrIdis+vF9H9PT3pfGqXvrMYTHBqLdhEiphnMKEu+Cek+eQwhp
2l/R1LiCPKPuLp5v+9ya2YN5xu3HPlUTQztYqRxiSU/PbRe8kUibfhMWNTP2gXZijUwKPJ1NPQrq
8LGYJqT9qDtj9iJhdg0ulME6thzLVUM93NO8ozpmWZdLBX7hWX3AnVyH9JeFrJHLeB/F3IFWiRR4
p9i3KcmINu5GGKBAe/BuM4aCiD04ZcRWPA6yPCvXU368WvKUSM8hntDEUm4iTZs12ctnJ6nH2xSL
pnsBFH329QHnpHMKnf45HeW0YfOCmXbrUl7u31oosfjWx23o8omNRNdpJ5ZsVHd1d+iI/J3WZY7V
qa5CdbbbLoCkCl2R6UioqFhXxypLB+xe6zvW58LPndlYmIuxs8YVfox2pLbN+F4dP6sCXnVHckxj
EzHQJ5aYezysPfN9kqJk8IYXBJIMPNJejUe6h3W/y82Sq4u0KnmmCaOaTh3nSnO1fcipW5QStDgZ
uhlRSEkmRNYRb0zcM7EgKh07feGmVld+67fyAlSx3xdHMRKX4hnS2pQ2W3GPhVj7wUa7QweXkrUq
T2fGzstjlEEVXjo6u0nlXQQ6xg0Za8Dq9Y+rwz59sPU0OumeK7i43Zfoi7fwuwAOgPs34ksSd0IP
AHVPwv5TAHOzrIR7ApJr5fHkR3W0IULjKY8RSx7Znu+jjKBM+zX6s3yn3gW7t270N/50aZbNDVKs
BC+FJdA+nsImljvhQLceBaiCEM8fsyMnnsLqqtigDuCG5cPj8fO185xQrqHFRnrvagxhw/b4sUqO
54+as1HLNn+8S2ArC5AQUjQxstwJy2+bZSWouo9AwrOvHvN+tsR5tNq8rjYbSwCWT8m/1qpR4EZX
yQiZDjma8RGhDVPGC3I3fchhuq66muOZxog8WYDaDp8ihv+Z2CAKFi4gaoSUlKmspHOGmH2V652r
8YkJEqQn+FGV8GmHjeEJMyerZtAwkscUOeO9P8HHCIL6ZkfkV+LfOLNB5leNvIn7iqwuK3AaU6vg
ctmUtWKzihzJK+vX2zNf0ymHDrcPeIlqaylc1zWTEcdQ/Cjg7TXlfUNlJD7xLUpUuvec7POKdUgt
FMIRiUInezRGinYU1k2wdhvA+YH7wzKmocEKgXpxghUIgZe6UuK3tBgTTXu32Uj0toiaT3S0kh2d
RzW9vwSybB43mpoie6xcYEgUXvMbE8xD0u7stnysZ9agJnaQrCawDlW1oqr1sWx/exWSpngVmqFI
wvRXqUbSmoStiCgleSkPEa9uRni2T/VjqW2c+O6uIIveXVxncVR/mVpgOBh+pT95enb1VI1a9vms
s5T91KGyiUHhw6HeaxtXyi8WkovZGOMHmrxbyD1jW1Aja1IfMcrPArXMx0nyEurHZ0Ej1W98cts4
TroxpU3VhQsz9pKWY43qTjrHlGs7mjkJOuAszTDtDgluoxkkuFF1ILyynYpibU6mHKNMQ5YyGoAS
8NNSCc3WZCtZudOuHvUt5Bg9s8HEsIhb41dzIxfCOYGJ7N2DHTx95/TOBWn/sFqMOIoBkqXStjFe
EFtyjBXcy3wLA0dzziozm23xep2h4WWGAyc3NUa6Ketx4QqCHJToyRnP2Zq7HNg5Rh6XoCAHVAkC
xwjYWzONjs7zQ5JP5+7OSEHA5Mf8m+wB29f8e0VtHljGYcC3TUwGYzU8Sd0Tg0dcqs3CC1fTB5OQ
49pzPThFCXrBKqa+gXscfUi1STJs6g+C4c/619Mrua9LaxLM2DBAY+lhI3yNpIK73CFoW91V7mw4
fpQqD+Lb1qslkyys//+gC2HHQo8e/SQ+FXOSs3C+ujzNK51BncSQ0Gtff9dJVZJSoqLdThQExY4l
sUXZcS3KMrcyqD3G9j7O3IpYPGl2BdJwbKQUCRPwXIvgcutdaKNmX+PpoXu9M6ikzbgZcwntkxtc
/iyiDReT/3U34AHvRjyylibKCROisLNiiFFQCbZmos2ZfSel9/pYLmafM5xf4rq+oJLhoQbiU/md
zbGFF6vhYhgaQ8GdaVq2JRwNhizW6JVl1tLny/1xkicgnKvEKWAVrTSForLxgkrpOQ/Sxq0/o7nE
4vLG/xUoQ60ZXA5t9ecttAQH2fKxFnmMPbfkbEk6bZJd1bu5+4nlesHHfk+XfGzcFeRrNdlMj8hE
PLAu/Wb6a5lhMeEoEM82gZSw/U548D2qwlX7R+9xmjbvEuVcKxqGrjw3l/eI56R0I6KhDbdZ+N1r
1n6mNeqFcd93ItpOTxqlCwgPWtAUh5SPB6/YGyC2XKFwVJhIBQBPunQApJyyP/B7+RydE/1e6g28
wSU7qk3UvHpnCs4lrA+EPGKGJhpHdsmKU1vty2UoNLERj5yEjRCq4iT2roa4kY+VRqHh8+b5u9Ee
0Mp1XWJ0dxVTe/LYk24T/hGoh6JWVVLvTfwzY3yNQo/z2BQrNW8Py2Oi7D9OkAB6Ene3GMeLgrRP
vB8pZ6uPsQHNcMlgfWC3/E7SGvn5VTd7jCaK0KRHzllBrawqg/6YsicI6QJrbYndP/Y8831RbJ2a
O0zgO0QbCLt4l8wMJCVy0lSadjT/3n8Vu12c8V4xWRc6hHS4KtnzIA+dCzzNSGLBM4xMKrfVz2gW
Kpwjv0t+KEsiPDl0ElyWfh9FMm0nv2E9DUEFrpHSUJ0v/AoTRno8ilmIB9Ue8Zsy4JIjGkZZI3Ss
yrXT3b0PvBxPJH/F+HA7qE9i5ZXS/wJbOu8I9CbJDkkxfHbMHWvi+DgFlgoWDshWbL26FmcO50Gc
VOLvOdQeU0KKaokiVCo+q9oZU3t20B7Vr00Awl4R34JtCo+cdxKbvVASCS2Iz/R75bghkVQ2GF3u
Ku/2EI0OZxUFK6AuzyrM9hOfqofwOBKf67KYNudOvVLsDZLr1j7acNvPOmmJipjd4+fvwJPn1agN
1S8YmbTeoKCsItfv1x3m9FskK5vnHwg+xvpYV8DQsKLGxvIApac3lREmgxUOdNSzGO2RdDKGtl4X
WJuygT55GnYawyO/kJhFflYSTpvQRHA/roXnFNgl0TucWTNnGVvVaCtyEKrGSxmJtr/DAq5t/65q
s5s3qxK6gA5Blw40JZYTSiGgcF0qrTvzGg9lyX3Fnj8o0SKkqZu3OLojsqVEBwUEQQfLOdr7Nrna
1/98DHJfivO5zUuShCIOJQC+E4HTPcYEGRhGrvjkm8FmjMFepS+pakid9f5r2W7Q+lMrOdEREyKu
f81DUbl+H6ezMetPcIWvDhbYUVoiHWcP+3creFrhR3O9YBAuTReLASf9qt1V6Q60Fnu/vu5TVIg4
Z4GdDsJJUjM4cMTQ6EapvREPjS1SI3EKDMFYA4+G1wKlBqrg+2i+LYI8C03WiiBqoXJXZZa444Nz
y2g7X9pGbGtBkGv/cnI2lEcY+nv5boDtuFBoXL+gkb66AVa4uTaN/uStcDTbQj9RRCpM1QI4CKhZ
ao87FwocZyc2EkF0bLB5BBsX6Qpb15jxIm2xSNP1XPlvvZ3fcOZZDWOQW+F5JcIoGa8iuhAX3XIr
CJj27sk04b9iSLjVN8qEB/yTVgS5yrnd2+XoAOiBRAnyM4YHcwsy9Du51iYV7HsJJjEle6Bds75k
/pnfMRH7ReEtnqY9GvjqHlEuF28OAE0wmGeU/HyXRVw/eSvOc3YBAEFCH1Z090htkXMQLXCIsqzf
BSUZ1NPCNxoTeOTUwpgSZeA21Mc7A3LIucIPf80L+hCQEd4fZ2ViYNBsf80l2oFvZRuNZSUHBbzd
kfRudZTGPlYu5X+tHSficw+rdgQOgH+V9Bhc7BQDSxRDON+rqM6tXDz2M9zVC0ZjiTUH1MoIoCdc
4g6IjMk6p9yOa6oCYqedqXntShQJmt2JOCAaKiGi5+9CWfV99LyrnFk4KQGa9G3hKxxO7G3XjY9+
2aOXDcxVJTkKxLeIjaMQhfGV2ctehiS8JpDs9O/KPMNCK1aBbwFbVsR2cSMD+jpYDW+aw0rr092d
MZtRYd3dd6KMFANcCvEkUZUW7EqgdjxIlWC0wPeF0+g3t6V+j6lG3367gXv6t5SOrMzVHGK0/Ri+
3K7jjP8t7KnOhQUBXC7csCQxDPP6ghx7G2HkOEGRUXlsjZF/ni0qca1pKKbgr9BN5LeVdM331TBF
uTpARAjW88TzHmB4jRgRwLvxzLIlsUL2iCthS7gVSpmNHzhF/KCLN9uZ/wjc8eDxNmWk6/Lj752U
KaufhIZGS88i0HSWbXdzXvDU/r2DjVkcBXD4gWineYiaqG4ZKdkvqw082kWAUjhjiUmguiTLh4GT
tQD1lApg9N2McTmSsUGL73XwrsRrDQD3+aYU/1vW6EGiOECVWwpKzYvcMrbXxkCuN23uPc69V5iB
HpPHKFJQximznsRJEAWn86eT8p2ykumweQoK9SqvhHoO3cIzOyG+bGpsFoNFwMqdKnOb/H4lT8Vh
HKe0Pg8jyr5b18srm6Fiece1mNvy7drUsE3dKnxrS/X17szrn5OpvRTqI0i6/gh+mJOxuCa7tuzC
TZd6buZkrAFw+7uU3z7Gtpa/YysNPm1vYktIZm8FgeAYwy9SXjyRTplYeICrTUKxJdUpWJh/yVxQ
7OwEXixJM5ezprSr+caJ4ruLALj912FdnxOLEnYCW9GylaiFDwSO7euBR0MncJ3WL3qLv1j+jQTS
7nBxH7PyHrMtcRpArBgwFcWl30wZXoMn+FlH15xAHht+N5XznWHh1dCcmwfEU3BnqT9eRvcpQWHk
j7la5V0px3EkyxQPFyv0odWKqhtlsVH65oMkbDcki6qv3GNaXqkc2hmszj6QQi01yv2blDh4TOw0
/AkfEtVShhWJGAOyTyQx80nS6Wx69CsEkGUM6ojoTjkvsYTToJGB4PADPjY6IWU0CCxkkofVYvie
YcoTESEYm8CghIC3cyqfoazDhQxAGSAtEjxoKgyGdz3XShfyRAroiq6pt7IdkH1LlAD4CGyG46UW
vi8OJo2yXiMFJ8fVuyNKk1mr1equaIl9E4UkQuQx63OIw8r404rfK7t1UO/JS6GIyqkno7SyEiw1
rn+Vhsv+myKceb1PSuWRG9evw1zqHRiuK5ievTTAj5nCTri9RAbKJ0wuwF4qaYFiIGUYmsrz0SXY
/JAnFrLlEGLnRQ+owNpybiyQhVVWFOSsHarhfBRD0dYbVkR7pF93QS/xnXoQxUGkPNMhujh6NN5/
MAkviqcYtZ0W3J0SHWpRf8M3+MkZd5pg6taBar19krq5YkMQUHA7iSx+yut4w1cidvmDdhlMAFUn
tNbZd0mljvoLY4fWHYVP+X1uca0VyIN/QEZ7kAxhhajiSrK9ONKOpfcea9tsj9HQY70npdOrcs3e
iTjvBjdeefFtlc/Oa5DijP3/j+pNHrgWTcJWG+jNR1hIGzEG0dkT9nhuCenasQztM676gWG10skn
fni37QKDGacTiKVVY+63olk+Tyc3zJYPmwjs6Vsjm9lYOU+6phR5UaeNOZJ+WiJdVT6h47c2omnJ
I4pOX7BFDo4R1mKtMsOhoVY5feD0GrujIsNt00611fnFtlxnahAKD/vi5eg9dTYuhjKPKDr5tZgg
LAXGgyWesNEhT11z3PufY2yrgtoEeVThfVqkKMis3YLZmhW1z82Sh5d7Bgeyk8DK1xvU1s3XLExt
T/vquzRiLmnc0l33fUMWXQWeyIVpNxRzshkTxlBZpsKKHbdpBsDcA6XimyMirWnue/ZypFbkL8F5
M87P7szXePTBWkxzXXf1XhG+yo9FH4FZkzxOsNcaCCMf1fwh0t6VAVUfS2RwbYHnDu7CtrlVsvC3
lzzXnNhS7GPyAREycH0rKvBXZYkADHNi7Kr4ehAabwPfsmfLk5Gi5HY5BnB7kOo7z6rhIoVGylPq
BabHt0+0jFoEChaezCOqDLKlC261q7wHovZooDjdjTvGDqWjr2s2hzMfxfwXnd6vCSue4DEJxyrB
XtcdyXb16nA55G4YqU03qdZRDRFkUN3G6tKGZzdwISxgKxnKZPrKUv/Yo+gqix/QAyAn+u7U4WvI
o/A/o6vb4+uqMTYF7EXPpkcqaFBiz4fkO9kINt9+qqau1xN1sPTvjNrMbJo2/70HBAYyh+IqBC/1
a4w7HlhKH9hp/xC46mPLyGz4xZ+hvizn45sg0dipAaFQ7NivoFCGVWLCGCWRvyoU6bo9OyoARCGe
tcGUS54RexyxXr689bQk4hy3Itbgq14Hm8ZFFFxr/3dOLrAfy1jnleRxqrMrxPLP/3gtlynpFjKw
mjAiwLhziigKo7j5zKty1X0rh+sXRQG3Zpe046oeP3HDZER/UuOIB2Qj+8BDxB09MFQ83u+gfNOF
ol974yEjT8JepPR25juj9+r8iF5MEHgTMBJgwryHf5fY7DdvH/g4oejuZ40SS7tz4WEIOjK4E16/
FGmxPjQXlwf2Wz6RlsvRuwzZ7psX3bpVueYkWj7hVk+kjbQSnxnfwDSNkGtXWqOnrr0hLPbVW3yM
tkwO/xlOZVcPWfb2w5Az3ZdNliCJGzcm5cUBgSBPjzR8xvV8nlQgojdS/yCv+jRS2eJTbX9UOamn
8C4A/tPuAcSA/PVe4fNViu542t8Xe/Cubq+G0CD2IBCM17D6ACuQpFrH6no2ZPoTOJcqShAmIdJI
x3dUCLQgTqZLRcoaj4uitZ0W/WRYc4OhUpOF8dtQl1W9MAxgjzqZM1Wh0WK4I+406eh2j8F53xWb
KtBxU6ihWjqjDeV56d2/3mP3T/av98gcCGQyBzHV3w1wr76Q+rZ00hhYI8kCRqvRcXHm3GCml8ZK
Y+nIfvLoZz+HXggABcj+yu0fkVxdIl8qBzbyESbRK8JsapdKsN5i80n6vkoEDkUMjbiL/rX5Oepq
3vwbPgWRyDjChjM1Wdc9Mw7wqK2tYZH/Mepcvck/ztAmKpaALNwKosw/KvCjSwdmdODCCbpsR9H+
CoTXlcMeUqj6vwzunbOrud2iAViDud7q6bBEBtbBriBTrW830YlFr6nJi7iVzstrNM5NkMZ3lTsy
+H2/KubQ3ineh2q93VDkTFElR7xLkpaSw6vc89yMC76cjyzCv3ji1mEX9gCBtxPcgR4aMwXCNPw/
hHg5gZknUCKgCXTTVOQkWQQFb1ZvaTBDhA+l5qrv8HKepAsioOvB5tTWXNqqK/pdhw1avDkpKt3g
9Q2rStPa2zR5tSHkXN/39QFHVcsqZPJokpi2grVAi2uTJ8hKiCjbpXBRyeBD9tYbvbhOOSWTHavB
dHNns4tbXHc6GlikroJAul3Hq+nsJuhY5a8QfprGSZ32W+s0RS6JjmqquRtxpgNiEWfi+wNAhtMb
NnEcCEGB7xGhtdYOm8URUfFsZXpppLgshV9rP9wiB7j+/g3ySZDrsMhf9r3Fj4Wmo3dJL/X67cq8
M6WJxMje4hu0akDP31EjfLoMUEG1aRmm3WgQzJojngkFxW1TMjRJItgbW2c1wLGbCAqTcngpMHHw
f6217whJKAf8IxSPC1YjOwgNzA4AIcBWZRxbK82uVvNQo7B99Bq5p/B+OGhvMR7K+XUFVaN0A0yq
8WD+AdHZP4LJ8tVa6mQL6THpd0Jy9Ul+xPKFWA3n7zZqY0sYFR7PXkD7SB9WqiKD6v/S9QUB6jEG
+tsYpukzDhmULNfUbwNFV1SEcZSvgT2eigG7GsK8jQuFmOrTAwD2nzwmxDjhnO4fhFK8brG4yPVr
eRTtXiBA1vyAmUnz5lTs8rrTg+gB7fAPsN9yCWlig5mAqfLHxlM8Aw2CgOiiYGjEqBGq6F/N6h94
1TYSkhOSJfBPMy5hjeaQFgeG0q1C/1FHr+MRCbauvxtxTOoly2iKgi16U4zGBftk6tHnnRToL3IQ
Uq1BSjqFB5TfTmekCFVY7YFedJg3MIVLgll6xmqKQNA8Wb63/NloRkNm3YFOq1OuSMy59DHrF3Z6
GylC727MsmfE68OOTRypMj6UuGocSbusuS5cMz5kSGR1tQ8VAuw96+SiEBnM0eyPeMR86Ky8S1BS
fQqZqJNhqELXCrMNu6fevzesWPU3YECF41ER+SQm69Eva3IdAD0YD0K+TtkpkvFiou9kXPoAj0B3
wa4NOkh+TCp0oGGFyWzHRU9+Xxt+RifmsBxBUDHBmoAlRrcJTXrw/MIKYIfxHC7rB9clSXhDePdS
1qkhEcYbQ3g9ANK6rRb43FsuLrNphBVPgS8aSrXQuk8HcMCiMhAA+OsMOKDyOTn3poILpxj2ufCx
SJbV+I21YSNm/kMj5w70fOMZBEpLbgwffaQpwz7gRQgbKTgSiM0uasTBqnwyuMxQKuKWKMN/Xd01
97TEHdfAL8t7xz/A7t/P1vE+IeyPgdJY+4iVOSBGfB9hgBkdlUuCuCq9YeHmOpzu5pkh4Lojd0B7
7xTnucdU3u/dnVecsChXbvzbRbIEcd8w8O+mAGu6b6QlAMNVuPjvmNtryEpZi6/kbOL3Xz6NY6da
SgPtJY00uKQTrHVyuO49wG7KNQEqN/9ICS9buzYlTXxwXSFAzYuPLwy6kDCLfuwLrimBWHi/5CMj
tqD+oBdgn+pNubo32274uk7dknZJsUK8P1r8tmfdrqgoitNqZ8Z5ApMAigXE/n+HMzrVQ03hqDwA
cKqX9reYQNP54XVcYXWYtvhFX4M7yh2H1o9SkDm5Tsye0gaZKIRIh4IaHukom0+dLDiby66JQsNK
gCIoJrd7s5Q+H6COja/mbH+sETBI6jK4lJC7aCUKifwKLEmLHWQz+J+skYm8/C5HkKXnMMxDvOE7
6mqLCgdBk/Ud8vxWTJ8sjq6qMt+dvoKqFwwc8gTPuYP5jhyyJgiGNy3UYPGEl3x2lSDtUQ9kLfM3
oKBr2H2krBDiL1K3kpRw8E4NUdbeiQnZ7Dns3Vrrij6e/2Xik5Ne6wJUeTzGWBFEHM1+J4/OrNJd
9lsPjzQjaE52n6yBBwfX/aLoM5EPAcVpWN6q4eeF1S+QPHDOoaEqGIeJozgJE4Lz0uo448Fc6Ht6
v45xpKqLdikQU9ru+LyoHT9ufYFX8TV8c1zEeuZEmi4jqY8RHK8TCKiJYGmgHCtKpI4hTWpzErM4
8jBpKXO4RqQvzSD+WtseDGnxcmF0Tsg9CV8kX/PGWBoxGw9NwkY7PW992fbyx22hSnAk5MVId8eW
fj3g+9rXH8g8fE0v5bXiOOElIeJznDt/Zc/xcB/oiAyZth905CB4BPjqiwwI3kbC0H69XMLa7WyU
yf4FGROCeMRwUJJnLYMwmDSqbwV1G8zZGYivsJc/qxhVTkiy6wwI0tPYzA7Iqs3AlHs6q/4R3sJq
Hx+ZRSsYmRhQ+SGxS/NAoARbLpk4LGsRrDwlfMJ7w678JBgDABncIHtdokGRUQGnXBmd+aFTzVP3
V+jb5OHXTdyHtomQmTNj8vXr9PI2yYaSrqORnNh3LFSWE2D47uVS3NsNygach17Rtg3mpmhZZyTy
nOmYLeoVDNftDuO08LSL+oUcpP+Ycit1/r+7kqpcWLb3sYdRZNRYXW7IHC59N8zUFNjKgMAqYuYB
cg6LmKKgPho3eoAeFe50EQa0l8HeDHzMg62jxrpg7YSF7VjkxzS8hTf0lCbXADrxrk+UmuoryaL6
YutON5N3ol2V04ZwB4LcnrPQNyuP61An8kCX0SPLDghH8xGK422zLtgRo2T3Sz+BD6tjT51x4ZKd
RdKSBwBTr1lAoZpMGX+0kLJaCpyE8t00XgsZ4l+zt3TMqdBo26uvr7NwhJGVsLCC45wxZ9V8OvYp
dVvfspmWdNDmccWhaNe318Xi/9ZAUOp3VzLtanOmceEeR5qQk/AUI30bK9C/4+jkOLf1B2pc8bvG
OlXesbTX3K4P0d9Je+yNVJf1tU9r3Knca26Lm9/XuZD4L40r61clGqdp3nKvg+Nngfhn/WCv1sAJ
YQnsOe47gWj6V0+9Zxj2WYxTL5EULRdFXXipwxsoQlGDnAsef0lpl+0gfBjGLHaHbyW0UqLmxM/2
CsQ9T5naHCz2Mkjjlwc94sPHQFlM3UdLJQFF70n5ZpHLi/1OwiQsXWXizP8ElAegzruVkI+JVpJ5
I0MI9Fm23IbVkphsSvfExirKotZtvsF1f6yfKz+0PBepm4GiD4dozMnYmDTsdO8EdmppniucU0qI
mjhncMOVT0wTxnDNTwFjNJ+Yv8cAsF4BrQKXElP3p2UzMuY7N9k5KMTVdtDdIJ+AD1Ux/wx3c+u7
RCc9Out3VNsJ7twyOCmb7k5JzgTc7/8gOX1kI1FKVkS5PQxDbfY8rsAv5fmtpMogOQkpOG3eu+uX
/UlspEbZYmE+Wayf8oEbbYGtK9eV3n44C9Zb7596gUDa5rnvZEBO3ORfKfcraHryf4lab4FUo1ET
/pn6OWfX5Owhka+rJTdYH0KE/Wg9q4ngV+HgBJLVyNRZ0jRyq7wtNsbP86V0cex9JmMR36HL6Y0i
tBZjnHQ9R4CpBoxq5RH38VMy/o/SRZVSnZcSt02VCn499FO7cqJT/esjW8hAao4ZZPLllSS4tLAb
qk7a5dT5sxDYOSQdM0lqJ8NoN5qep5dgjIuX+DY9m5xFNybGqejPUc1pFOZxsyxec/eODH0e8cE6
wxiDv37IFSy24Bi+4c+bpGPM59jEknen9xGxW2c0Cjace0A0kmuaVhaxkhwCqAFol6Ln6koweOey
gaQlUO4RNw4ma6yaleHa6h12VD9o6tJUdhFJCUTKn4SVabkx51Spr4J6Ioggti9dkhXIFbhsOahn
Nk0pNM5unVXDQ7gbLF4BrP5Eg+HLM3a7EQr+RjKWwBZIZvtXYrTfCIQzxU1Gy7M0V/OlTjuTREQ1
Oi7xOGJRcei3jJNlLHGI0HU51KqvK9QYCpUVvPwjYwHYvUlYE7WCkcan0AYrgk+UfZ9v0Rcia1UT
Wd7YZ3sTAQ4ZvPXRGY5BODgvz87RWuvMGrDvqs5WyvvUaC6k84Ex2VyJcENhkA6zFd3OE4lyrU2T
ryfCF+drcC6A/04A3nFU1nzh0eFdxLblSBkefd/hX6TELZx7jBI0HcqYBIdhxh4GAvIK/8m3kFld
J7Vs9ZZ/fBeKU1APRxq/ouYkrvN8MMUXKIulR/jhUtP0h4Di6jX3TqZhWSjnVri+D/xoqa+05+90
yC0ewa0kW8l2UEUNFhe59AksOE6xebE23ouP9zeAYtIxvBABBPd2Le3y785NZErEuOdFqRcfcHou
IbHpaf8qgC+HbTuKgQPYDDKZme3k0vLdpLb8tDyImtPycVF8BoqheuBP0WxvBPNhcMMlhxfKu5dK
pyqf2iuuE4CdjtWSsybnXItxlPsyhMZ7x0TXKfqTzUitXKnWmBBSOFl9WWNmx9aVXCVOhm9uwiNH
rnKR103C2DiA3yVYmfocTIEYG7GIhycV6FXTHTXHvl5aYRPIgx7Y6dcOUY2lYLV2r20D9vIrkKpw
K+tCcDrKsjt0KuQQe1JhbDBMaRV8Q+ZD2EHbokVg70gJdmYa7CMgQAWlXQbs7TKyiXcRX7yT6uYZ
8oAx08Xr3ldSmTbggLHvb/4muUQNGUEXOFmnthCtUtcIrm+UVEZIJat49Igoth9CG6POAdHp0yM9
Hf8DeQGpueKnEmYqJvwuwsctS7ua3rijN4rTS1d+R3L/hvox6ipKtIjyifV7musnMzID90lwJb0/
IJzbZCMZRE9LGmk4h3f6mMGTrlVrKLPaFW0ibe3amXECM99kunW8XJ6MYc5BeFoSAntJWw46MaHq
nbgQlfmQgCkD1P91RNOQyW0kWGRn2kHka1IrfBfe6Q2XkUM+LChboQRmsGQ2m7bpci9rZrYWpWeZ
4RLyFUc3KqcN6J/OS/DdRrXwjTtrCIK3r2wnCwEma8mVNBJxarFw2M0Vgt4BdAPxKlDJpF9wcddW
smPAmDgmVprdhYHkTIpTy3QxreDVLNEEaglSieMf8KfKRgN2K/WkSOBLZ5PvAo9fVnbSmAWgRmIz
yYDWnhfI8xniRI3a4mMhcFoyYgEh6f4+la3o5oyAuts7mH2d1HWk+7RPc1rOBnhVjk3hoqep26vj
53o0bRArRyevyQQOmAbiTRh5dvQ1ryuxy7jb+tLOuuYKssXmZJYohoyrjK6EKjkn1H6Mz7n9kXjT
jBWf4E23xe+ssnc3nt6tiQTa52DI21FRHwcIogQin5Ue/sFmTCLbODaH0KfAjndnIue8DM1ZXd1w
p5phOkgqwdG5RL0kmu+MkxYIjYOHSYxpmFb0d/OA5b1gUZIj/xw6FvUiWsXl575KnsCRgDwS8K9S
xoS6xXsuuQebtOHJ9CnjCi/G2Lt7Ldgo+dl40EWpY5fgrfrXeqPsM87KV/9s8KDwnb06oIqdtPvT
XbSIm4D7V0rYHVQvYhwht/hOCuzzZ4Lj1oIkuGXxhech8PQaNI3+WXvNKeBm7kq/XKoZsgGnRzO4
9JEx5d52Ot+qeJ4OL8149yqQhJO8rwpTeTFJDlBRLKpxQgBfK491ZBkmpSJ85vK9swYooGcaGgKc
NXcvehEIEbHzM06g72P6ojkKJYe1fKV09HyVLmxqg+W4SpOn9+hjQr+O183FIvQPy0cpJ4tzcO6t
QsCmCJP5PWU/a5xszaYaeJXSWwx84zDzNaiA1NojN8gCVoIHnUDfBgS4nKTpAiK+3Ly5O5+1mvBY
xQlGTGEE9t2d0KumUucCh6BOc0EB0Y+wHMVB3pjz31vPCVWKEcSNtaLiaTwf8NyJUNdNOWrUXzTY
97BMA8n5MbIEgk314exL2FC+I34nbpWN9ZJKbZpcgWjWDIeznefemjzz+vILIQe44FpqRnITDE5J
y7COkWN4Bp7zG+UOuAhYMk5gvNzuCNSsDRoKQb7T+DYP07x2NMBUMLa/6XnsVo4qDy4vUnPFnSG8
noNQ55Y5O/vu9lhOVDZbwiD+ym317PjRP/h2OUn2mmJuZb2eeOjWfbe3wbiWtM1iA6g4ZcOtl7Yq
jqbdEYxW9ACoerbGNA/2D3+0cyCQC90eBz6k6f/BaGWQeba4qD7tCgeUsdXH8jzd5SnZz7m6FgSt
/2QemuCOQrK4vPaC68QhB3GbBf2iJx7hgYNjWZzjnqAbtHFZHW/2pPqp1EasBhuLs9WmFSZznQei
Dl2sAvnimw/SQl9N/b1kKRH/gvPOs7k+VUQUemnJJP5Lk813Fx/KrvX8WIknuVmRBBIXT4tQW/pz
cKv4sBU3OfV9dqQSOkSsR1qGddGYlX0gbyo/NC/gsE8Z7v7kJiGUSeJ0L45UQtOLqwH+flG7VQcm
lsA56NaAawrjAabQnGNm6dgTmjevqlcu7KxWF94Fu7DjRBf9xbt2qvwtUkSdRW22HIvxwNWFXXyW
0Vb5TpgGYpD3/mYlrtfsV6ELet9jnVZPbEwo50ouNE1eKLItHtXnSmXCsp/NDvacuOEUCWnBtH/3
IYwH6TGCmna4wXJmE8DaJUjsh765Lto0KaNVd5PR0T1SEE4ER0JuuuV4ZXDLgV12g8ATcf/hX5RV
UhAsQhm7ThXvKy06rXIl36/XGgsVHKMQQ6WrGzyhKNt5+eiOTbEsqote+ruGk1ZClmNxhrxx7aQa
WTlO7l6vg+9ZHdzOvYBIlRx0EBF35k2KNXCjRDRTOw6t0dRiDwqSuLxIdS1eBY8CgMZYDlfwvfLP
agDV6nfKrcEPiKfhI+W0+9OWk1JkfxCS06BibudPX1u6Yn7/CLaB9X1hAyUXhc+LvutcwlDH1ew8
en43FADYSNNBgK/Vl/RK4v1qDgk6lTQA3elP8vGe1yoy1NrYrdfRs5fskgNgIi457uIvFf34MD4P
vflUKcWh1NZbprdfjF+wnTJfIqdvMkFOYEn4iTEUuJZYOBk9G4P4Uzj3nTyJzfNPHcltyLzhl2bn
tY2tOO8W3b8YvfMALYx54Dn+xgKaQ6Y6Docinjmlv4GBroqjl5J3lmImLfkuU+gmbZeNCu7/NZom
FAcn2hVGGyYQ19S0Kacly/qw6Qtc9G2KSkqyviAUIECKkAv4xrdQiae0nAntWu/2pR6/BRzbd4ig
4R2FgTLiLS0s+qxTunuWm6DeMRV/3OCNKWALEDq3Di3kHRzG+91VDv6GzJmibm3jlTspbQiCcV+8
kvCeaxlUxPqpf+zPs4FFD4KkZq9MWHgbIwmkA3B2qMAKZUN3gfOME4viNx5ngp5/8LC7yoj0dTL8
ESEqYHJtW08lA1uez6qzUnb+sXzoWE7QQdEYtgt+EyfxBYrM3T7eY1k33myicEWKTSRhffex8men
4OAA2cySkcrfwyjcp8ohN0QUYrsGn/OtCQG0V/LGeD5pwsFoAff1K5H0iDR0EzrUnsGg0dTDHzyz
ZWfAa6VBohGfL2uRxr5XorqNg/Wez5axLkLr0A+OZ7HAhG5/j501Urlp3dGym5+tG2vhsKkYChY8
uaBjT8nWqMZ8YzuvjSpjiio+6lDyDAya8d/ZQAQupvNKtL5hDOJjVIppkvB0bt8PGl0UuUTdAjP+
YJSXDwfyNe9ooNbrUBfVB/mZtNbn+Ul7T1KdFfdM2y9vbMTZKS9mSxgqBFS2LKb1Roh3ea+IRvNt
lAmOwm6A8Xl8MUyobK0V0zQ48Bpx+ICLbtDLjFG0J5Sh8alswi7pjIXHuf0GTOvPlXp0p3ieVsdT
XWPUY/LyanhEvvGSAU0Lz5Kr3mg9TJLFNHXUh6kACtKVKPZ1LuaZptba38zfghTEDoY8ilTcdH69
0r8MwXU5CfXkq7qiAViIAz9KAiI0xH1IOrzV8z3osqjBrGtOwKlPfL2U71IYcVrOg+SYI3WiD+pG
XrVtj1iLaWEQTbgdCUcddeT/KwZk1eGUgFvms7SktIj0L2/84mnjIBV9FRvdywdtBc6juGdV6U3V
blVhJDmu+gVIHzhNT9wb8yuA5IC5EB5xjyFHyfjNuSmel85lQHUwiv2vqIcb24hE3+DrUG4fwwP1
XfKaSqudyBFs2hceh0K/2mmR+DobM5v4E2zdlfYpjbwynyiV7umSep/0SuBZZNYwOElA3dNlOP5J
pVN0rgQypI+oQ9+JGieVNYustcydS5FVbE2cRRkfp50woURxkJ8c5BMsIxB2PAX9UByGWFmwtwuQ
LinDKbTTYoMKZDdU6njyfDuDcD0rpEaNYX3n2jNOcbMnuvLcEZK+KLJ8gq3lUXal0Fmmqz4yqlIO
p4nQ0kXhA7jgvhdgOtUWReDFth4r8sndERxMXGtq1RqAZ+zDSbYQCaHdMapb7iy7/GHZ3G2hwb69
vfDf7QR0lYlFf1c2jxEv9n2vtNkxyeTHGibGpavTHOI6MLG8axFgWOE8NmMx0XeLy+DOZuvOUrX6
+UPYvyNmWGh7E/OANn0ivHj58tPwcvvyDtpo42GqbiLRYynN88c8SnRPHNSHLARST26/ixSlkdt+
3fQoGdkWmrEsrh+GFr3KUxroML+Dz+/uAy5EbAkDprfkSCxnXYdpB+JSaMv5YApVETCLiv1qZUrs
F7v53oOWb8vuoji9hIaEA/F4OJE7E++0tXOCUZASTA0j4A2hGfuo9BKudvhsOvgIAqUKmd9TuiHF
sB3ywvbokmOYpIA2WTLnkprx94waynvzqy3ekdH/w/6EhK6KMi7A1GlumDYCMGu2X9ioFMgM6uMu
gb9xkOmF2dPkLuEBdi/vSGfbYyvVZEt/X0gFBZyL+dNBz/s3x34rc7hy9q1N+7gxSVd/AJ9CIart
xTAPvUixQF6d2YlLljWCl6+mD2f6Bbjm4yr85aYWSTghPLlTkCFpHQjeV+/QzDfYa4MyjHunKn43
beM4L2VQoVwOX+2WK7JhCZjdwBeJQk4iwA3TBM2iatPVtxiNrJYqt8rdHNSwED6vQHH4uHpECjeY
xhg4qvnvSm549nmi+2jgces4QbSEN10Rw6J22kmz5qzwDeT4bzLdRu6/owcfnbjK4SU8i6xLXJ+V
OAO43mGIHyUfRJr5CzJO/9xPJ1AWcPBxM47XD/R9LgzpmLAi+gQCA5Ohf99UfGfN5Okxm+njhwkc
gl1LPxGFmPlnRJIT9CaTxiL32Mx1xvrOuY8lckTIuQdd3xKraXWHCQfrkOluwh1evTwZi8XPuO1T
rMHCW5tctcJAyPcL8bWNGJvQw8C/rAHC2tClRelYWULJhfMjvu6eYv+9e35hvpdJenThPgiM8SsE
BnJ9o+wf6cynVZbhBveqSG9BjQOecY1+rG3RAl7QJYRUAGgkB8qff57qZ8crKw6SOIaB2imfnvZo
+rEtOwZg8y3KkyEGv0L6hhdu9cNKlZHqOhP1GKw6NUehwHsV5a0HD7vsNHoWJFVwxAEutglZinhc
KPhQ/0O6CxxiRuSXzm4EnGV3pRK/imIn9yBbJja3PNG3tk/0CplPfnhKx1i+WL/nOcIEg3juLSxm
bQ/BeqGaRrRTT+ekQvMD6FXgnp3Frt4m8A9cz8EQW8Hg3O0gP9RJiuqlujEUQsY+pezHOemx5MJ7
hkd2mNSNYso5jqGv7xzCT4Q4FOAvdKVjL3QtKuvLGPkXpFpEF4KYvgaol1VGUFPeKADcKSVXMJH+
eD6qEL34bA77uoCh/IAcdXV+pxHXJMmV86CjcxmSsy4e209b3VptMOjymVtBMOB2+Dea2e/4/Ot7
93VlE9zZjfIKVuZPuwGixiJQCxLsMsOBw8s0p3KYB6Q3yPe8TB4jxCKbRze57OHP6avAVbPHwWwY
+EeZVXmQqIBbLEpYnSX2I8vHnsylMPcaB6iGGznf/f0ORoNDmxQ3A8HiV56qpjSJInNVWrYkN7XY
8UnNSNGMcpfnnBnTKYUYpJFVxbDqQ1EJay9pFCVzqV+rQBLhSxJ543tGPywiHIpyHT4r+ljQHOCP
B7S2bNoMUjHWLaInWHm/YhLrBw6Q4WlYN8bkN5WPyib8Tdg2lhFxoR+vm9cZa7EErwFYfNNwS3eT
rYoKkP70zR1k7pqqKd7JuJ7WfdtkSgAKCCoE9c2Hmg7ZneTiViICIWRTmxxgIJwLIHuxbB45ULPr
eTpXFFoicW16BtuI9nx0YvFlTy7Wzv3y1pbDuP/InRgQ7Iq3muhvjpOW5KNnBEbHT219/tV/ha30
SUXX8KYKoHrgP6T7wPb2Knt6FvSXdFaq8jPbCiHngH2lIc0dAGivKct4zZkGJmODJTBPruGd1udc
IzT12Sfhf+ev1JZke2dRk3xP1C+aga8fiHB43UOa7cq+H0kDWbgjFtmusnIx3ITE6TMpEMFNc6nG
A+/1E0/rAa8HWmnX7wmNJQD4tDNqiqC3TXQ9kl6r/+1Bbjl6Lw4O4XrZ+4vJ+uKKNQakythCZTSL
k9SUkCaMuu1UyB3T7efF6XC26ZNltE9xx21bD0muOEccrlKvkuL8jVq91ajGcaASNZSwf9k3leRX
bO4zzdv8Xnpki3ryKX5rKVUt4MdWsxJwlruaO2XIRDUrf2HDtgY1dpeMZPW6nt8B4EIyMmJl/i1r
KYmyyK/jzcsWxrnj9fKInLDJKMJm9Mh7dmedVmUjFiR/fPsnTxCwg3g3gGO3s77HNhdPKPKhGcop
FjyQuOtI3zcVcoFhaAY2W7+pCg4BiHNz6CTqh73/+PEVWj2R1aoi53KcobX1rFhL4ZJXfWvhmL7a
VfvqWe979OI/JHRfF1uXRmeLUWDQLKRR8aDiWWZlUAFh43cGyZ4VE9Y6/t1Vb5sMhe4Z8WSVZNHA
EIi0XdiCIuDUGfyiZPLm0+9IonWqg0Va3xU2uGsf96wKq+mul4U9GSig4wtugMrKZnJg2xpdpg9S
AiUKQY5NyxO4F+5X4x/z5XF0xgsoMrsHHLwjvuxiA1gDebOBHgRK8QrCpdbOvop8qMf7M8yltp+r
NmLyQYVJrLtxlROrLDiaCPGwx/ePvAI1YzCdjdrmGrTUeDgbCZcO1cSD0qBcQhyCN43GzuniT/sm
6O0uy38Gy8j/ZJ4YLl+ybAzBKcAi902gSxqFl4jTlRvEPtBTm9BzOKz11OPpEOU0BMA3qw1iauc3
z6Jn0XXMjkkHuiS7n/sOFH6k+KdwNyQY5s6Jqm0QHqJkmPIGJDhuG6wYVyOMClSlJyA/ic6gyykP
LPVT7nNMLRCiDBRPctdcy1oZ9JPgr8T68SaO2f+p2OWSYmTeX/yePSZCWF4LFYc9ZxsUGetZI6RN
2Zq1/4kppci0zmOSDUImmn8SKSMMqbdAufIKQdQDx8t4zpwnbOgSKQU17d9U1HIVMe2OhryLDI59
ubmHuUpOsMNdLdt/Rb64noE5HENYeSNZIEfY4lcCxwGjoGTeHJJa01y6ZqufpS21vllGUa4oJjr6
Dh8p0EMAzvmlZWv0l++qWLD4uARGf7wMCGq4lYw03jBdHXNv+XN/3tpuIongC35qVx77DA7KNBFE
YvQq75cjpewqIchwC381s+dfWzdE0i2mhRmrRsWMS1VdQS9HOSzVdjlCbX8zSRdzUVghqihO/JME
moC6zie0m1sS4X6GHgz3yTlClYyzIgdP107mG8xOuUzy07uxeGogroqMavnzN5dDqkOdJ8qB4+fC
whaXVw/6U40P/AgsZJQeSqbu4cXNJi2pq23EwQrns1vKpcYeraz1JQUJhF845QBLJREaTTS2PWLm
JAZsFVnKBDLe3muhkm1YUqoXJbExEGDPo4UQg07rtyRyP9LmIhdjupLojjZLnZyIAhlx6V9sA5qB
eUHHoWU15xSR5D2tI5q1QHCdjuhnqy+mYdlY19fNOPTsKo3qRtKQX/E6P610xWponzfnEUkvUSRb
lIJsy5qiqvhG4bp2QQTGJNLher+eiOqxhcZ1BlynVaY06HfIZKdzE8JOiTMcXClVLonevD+XMnkN
e69oWmZ0uC04+oMkidYVs4C34hhrb5H0O0H7qreQuGrUHuz9+DnEhmzs5vXvJsza7SPrA4CjbnyX
gGWtUP+WL/cf2Uh9LngbUqDac3ZkzEmuVKpYnFoIANA/37RfpL8LYxjrJHupFOqozpH/ltERyugd
GFxQt6Ay/DKRa7IHzKVQbwpHMC+GShSNDr5ar6Up/wTKPqfHlsNXIXH9bqG/NfSqsVceDBAoNmAB
iV4k5UpPWdJ0Lp7MvXUIQbtZ6y+ZZXAt3Q1LmPgPL5Tddub1zzCea/tk55nBOMbZnGPN7wLqgxdQ
VtA/XP6HeNTtlbnr9sl4231r+NaOQE2OGJDY9nrHbqVvulFNDImMqpYtQMBPfDXna2jqwwE5OXoV
Uia40eoNJpge9LXwAJnF0a/PgFMh5mUYZPpSLJ50hMHX0IX3ScspSLl4codSr51rgZMCNEhRjoKY
dRnmCMD7zqziZDTsWdZGYKpNbbzhaS3EIGKl9tIQGR20xAR97xo8zO+MpJi/HGmfnOno+m3ugtw/
Jwi/Fsui2+12SlIyNJmv16whnQsi97/OwfXoQhlzx6vmmCEeoToVG5fEyN3tnFZ1Dkv+TFtSABR1
5te8PprdJPJQEJbNvYEAqhq55TfDtZ9GuXeBpliDBcaP6rp1kzz+Jd/GhEv+8IcxhW9OgnvgpXRW
75cUVWLbSW7OKhrwxyKeivrgNCe9pWMt/YVDWmkdHoukqUeTXfqbmmwCQ5Mnkl2mo/+3i2o/ArI1
xoVlJZm9KmK+vQlb9TwNZFvVkM7mNe6Mp4uNO/7KhIM0GA+8ZqE/dKIeBqBuhc+s0GLsA0AFlh70
LzHKOPjIktVp/yAb+iTpUKLnAxKM/fXFierBFAv4KM8S32Rww8n19DIiybxVAe42A9Kgw97R0T7f
GMU/gkTmoUOmT7kQ9aRd40t4LpFXkf4B0lXqemiPOUd4u7UEjPtU+i4++agnWLbcnMgLBe+BtsYd
GNT2oLJ0oCscYB6vRVmTcGAWSZkk4SyWF98bEwDss1aRlCC9n+A+N1qjcIPUqbAkPEEPg9hK1bbN
hSn2Z+M9I4XLCaM1qkS/CDS1sX2wZAFAGHUyUU5DTzInASwH9XyAcp7gw4KLa6oqCnMLGwEpkiIS
GExhbvgomn99ptPDzXjzY+F3Q8YaxGma0CzYfxpwTx5NzyMqX4h0+ixUAixTmhGqtGxR68V4P0tZ
Sph3dqAicP3o6EksE0NgTv7EalMWu1gIAoINC23ghfaNcwRL4Hd+F2fdAVj01DqlMgavN+motm+U
2rVMpVhUeULSeRHuVHDDbgu43/Yhb1qh06T7RFWKJkdGBU56AohPqoBDm3/bmVoUZ34hY7+viHer
EqBQRRxgkgj0zh+i2/8LjGUBy1OBxjFTRuqJDO90VnZmYoGCd62xTAcgE5cKd9yW4nDO4HNMlnLc
xkTQ07YXLKCMrv/nlyKrO6uq+M92VQ7cRgB2PAtuNzJE1cK+0PEIfmsPJM/bPvMIrt2GmQbCDt/s
eQQfYrQntzHzjuaxcTAIoHkB6Q4FM24SCWEMV5TIKVRVRsflHMqvqa2Is8btXe+zXICYJbhd88k1
5n83ZbNUvzjwyRr4gMy51iZp2G++vE0/xrQOtkkKEGeMgWmKu0cnO/xkFXwveaT5+TPTr7KjU/SU
L0FTGmnIoEtXN+dxtYll4GhiY/xKagAtmpyrnUyd3c8N/Tl3yM3RdGIcQy6ys6rH5EHL93W4s17T
XNIPk2r3Cut5KYIdXdB1519XAvAkpy1YtQMAoxggqvqgfhOhqvx6pS2KUE7Um/5JHwcmoc2k/fCo
aD9r1MIWm69BRfUeiBo+Zg2d/gbTZfSG7DtUslOZTWleoAxKZPNbr9Q1YpS+jwxoO3QGCHDjpXpL
KQyb7QNYk2vaTh0KT4Z+SFLB7tBGOiAogNofS2KK+o6ZWWopH9FRVvN2A8LsU2dn0eNsU/CeJvOn
I4Xn8UPdGqPXFLZ3P8xL4eqcQR+4CZQsLGWGaVUWKUiIDctJZFWUbGfX3BwhWAaMP2LwKPO9EjHR
a9pgZFn+AXS3SItSXPCTDduP7C/SVsMkTVL5B0e25w7OT3jHNmCBpKfBTaLZ0SAa3/ZujmAGo7y4
hfFxVlTAcurOoFURN/z5uY/uiXBv4pJRCRvAkvHPaX9gbsCmhA9Z2OEDp7bM5WhDPN712Tt2rA82
hSDUfLNDL3b9xRaHW8mYptjVqu/3CoaFN9CMEhHufq9VkZY2lHd/9Mdml+BSIIqrznvARpoVRebz
tcaxBTsTjMNQXZVYiKy0a2+ry14vam2Crtl2o6SIC7ODcPpuNfKJI+j9JXod2/k8CE+nFxP8yuXp
b0hIZxZSlAfJvyDrggMAIZ1E1ecR1wYInWbqKKf9lzIkFFaTqh/TqUQYMPBo7NufQyu/iBjis2v1
fOuxYGujul8Vtr/3HeT7pjuVL6cGsQbBw9/j3tTqRzR6jhCvmWyPBinmiFPJUb0px4b6U1T7zxdN
Yhip3PHcaE4V8e57gqeIQ3w1RS3W1MmLrftad5QRzmSdf4mim2H669qqkQTJocIiTaFgkSFs0tAX
i3Wl/AcLg8nnqaf0LMLsrauAteo4AUGOGtRC9JAg8m1PFe7miY81U+lGUsPTPFX5OECeYNjUp6aW
lkldTriwD7kQrFLAY+ud5ONS1I1n52S4ZktT8YPelKWvoFxwnnWoIjSKpdXP741QjaOBkiGta1sV
sGG4ka69OsMjs5LRU5jvpa2Vyql7ioNskSzzVMzRKuVX86RbRTTbLyUqCB40A0ISKgraPLMhwdl/
p0HO8VrIGNmBGcPcm1az91SL7S/dD714YQJqLc+u3UUZpe+b1AaSTkYCb7M6YPx3XBdhoSkobttI
Jtd5WM6YwDmI44K7ryt6WJzh+aelOQdmaMGXDwvFSXhLr7wNwy+202mxcx1uECVJfDH6bLbzW2WU
s3IQ3mADVJHke/LF9ZyBv/Ce5Go1gEmlRcjdjqclXpG7QfTE3srsyBH5IKnXwVZ6ZEJ33DiuuP2a
b0arRaMpTSk95+9z+M+s+Afuy2Q4S+8v7+oJuvZNzNEVZL7G7cSMv7B0n9XicgYJdcHAMbUssUpy
ZW2CSDuf9b5EJThiS/T3tfOSLYbq1JAx1+Klq3azQJHGmluuUcvK2Ms+P/t94OVSTDWW88xjwE6s
sNmXEPey/UhTTNAKGHoJlXiXaEKmsIC8c0mK/VoKN492NEY2ENSHHY5we3BuO1RjIjx+O4Ns+8Eu
qmFiTB3xI49t1UfjREb+DT+WaMcABDh5TqdzD/QpvQi+OinOqgQh9+ccKhrRdeoG/uxR40XK7+xg
UhutoPm1+VWh0Nt0kpidQTdebeFDbx12RGGqXVCxRt+btKwTfTJHVLIgvOn3uw3q3NMhOoQJ12NU
2CQ5QV8QX5n5DxZG0w1H7AVKvfdn/mj9rw5wPyJbXp46eRQoNIBJRfnW8zCk5NpsWXg5TXlZv0F1
kwuaUoi/+teklJWGGr+6WEukC80TER9erctZieDC2npAhfGr1GSiY4/zdHOD6r/9Dg8OxUfd51Cj
FbNduCGw5iZAV9jP7bi9WLyiAdCq7+PSDwzUUd92bbTxhqj+l2MPkdDL1BsEhk0TH2aJA7R82ahC
W5jUvx/1eT8ttwO8f/ocr06LkBVeHG3GbtBMVfzqDF3FHAuYNHbyOXT4+ya9/Zq8CMAi4s5SXL9l
tMswF+eMyv7VE1EI37fSzU3bLDV+VdMuMH3NLF/tgRr1zU3e8Oel3XPJrqT6nMezgC5YkqpcAFV9
5mUwOM+C0GS4fzvQS/0zbpF4IgM6I2SFBmeXm57ODOxL0QnOH16c4vo3izoRoh6JoOr/08/67qDs
BLCftVM2jO34DF2mHvDNMxXS7QUnUTydHxfqQsei5yZmODS7NsJ5DRlmbEZ97ed7FNKab9Eq4fTY
vjPZPEg7U1NT3+k95XEVCrnYzI5jrCs26ELW1nbq7/W19MGzgh1YDL4FpBid8Pvq4sunBP0S456Y
iKcW+n2jbBdgjswqCSoTKdxK+7DXw/IUhFPBYnunYPBnzObyDvkU20sm2wjk5z3NxLoBwxznyQZF
CO85V7XFFSJJ2qfIyf5IPQ4R2gnXkvohv6BYf4RbM1hhf97rDSA6Debs6B8im37y3Kra7QYuvim2
V8z5HaDSF/kVvsXv3Xh7qQyD0JPzgLN+9FkGr4ei96B4ipZZ7cfAaSombIvjkX3WfnZUxE47pHZL
pHesPgFcMG1WrnoR/g/ISDqV8eTT6Vtfwr1KvBfDesgFxiCRsxT5KE2UeqZgl8oSi7rIW+gifKDR
i2pPX/FxFGJj3J08ap7Xv2jO9ldO1nxqdDUKQ83xq84S3d2MeJ/JZpjY8L9HB1+aSX8WsKkoTXJK
MUwvWPeaSHrTXNJRafT9BiSjI2YoRqQtCPRFU1PIpOniempbZT6xGwdqmvxmSu/uny9hwAP3SDEy
w3lmc0/CJhJGkG8yKcJMXdhlS3I7swcm9tQPrlN8peJMddUv+OTWTYxUX7sF7FwnV5QOdMkSFp1M
krKiP9J0jio2ku5nZ+DG8LdM5ilKCcrN2b7NjAmClx/4b2JFNw/RjhB4szYj1NeE3yUWcZu7+bwV
39R7GruPc+DMqfKxNaWr3Xxjmc2YVGkvQlBh77lRaml9iWXsQGkqkUtMPjuUn9XVbtDTlGSPB9zx
I5zixT6b9kV/K5/iKsrf5Pb/LRWaMlOMo0uN293F6TFUeMN7likYnveclLLNif7e3y0o0wbhVWWP
gd9CIPP4Bt8KqkPCrK6r5wpZfUv8eyR2mnJP4yl24qD8NPkez5ZM1qPJrhk/Yljw+jVBunnw2wmv
bTJF+iMK1+NPtLXw3+DegF6y/6SqkIuup/T78iCjGafCXeJHlEV7fSONcCyWUEec4rHBUvPvzv5t
OJ1JO4LRiQwoTldWrIrkDezbazFwOSX7wqJInlwLuFdVnu5LXRF9Iw19RtFKHLkCfDRQv+r1Rkuk
ukhIbBzqe6nhwTx4ThGUZcHxb7oF6nPrMyAa1zmBaOF1wFvPH3jpggSsKe1DtwTPsdCfkYBSq1NZ
+eAK0sXAemGcUu60HazZTDtBb7ZcAeXUH8YXHhIuWKIEJKXahh+21TqyugJUEYUq+kR8ZAvYPFEU
Afn/h6zr3geUaSP+GMR5Cv3F79pQZF/eb5a1wJcFD9V9JuMXeAS6IWx8zmgsJ8hHBLTPNbqNlNnI
Iyx5d71V5nOkYbiIwDfdkMwTl/2Xn9AQmv/sKu9vNbBiLvczEKRBh+ElFDo0HDDLZblui+9enCnu
B9F7wcB6nkjapKJXxC7f7r3lCcsA0RG/OozEDcoGxsntVEzF2ulrKzeu4FRlZ4YfsP/jiXlrFc2V
zYlyejU3cmuLa1XackLN3lz1UiIlIxIhzXyY40yz8RHZ16jYn6OTvf2cRwjccB9onOOTo2kvuiX1
EA7kjxqUrz5iHkIwx9Pbu8E25fRkI27XZHsdnBZRFBm3a5fN+afzF1iD7lYvyWe4wDFQAGhsVQyk
w4s3Dmu1c3lPLh6q9b7HR3KS9Vjth9WRWMkxKXK6y74m/FLDG6n4ttM/AiWGiz7GZkNFyRdVm+Kt
RC57JrfjaqwIZc3NVU5ZfE1E7TI8/zA63MIqBYyg9fLpTsXA7208B8Sgzg46r+JoKzwF8xO1GK3I
YaI1BeWneSnl/aqnMzq6Ko9NsKt4e2B211fqfN4qR1WYwRzKaqUj+/ydQi2AtPBbmX7e1YA8/CyD
FjN9Za0nGuRbByFhVNSnRhhSxs3bgv8Ka9ay63+LPJZYlEW/FnCIGUsnCJEgsjExZHOuuGLBtg3X
pUS+tz2lxp2WcQ5RXMEn6yQIBgj/Ubi8+CSO+IDKNTt4HTzFMMD5fnMMd0b86lo9W3SoHEntUyk3
atAHsaK3YmzPPcPmC4GE7B/y+XuPBlJgIvNF4jLzp58nJsbbve2GZS70kig3FNfC0m0vfnPNxari
d675Q/IviDWFZ8B8wfH5e4zVrbs+jJXjPGMdkY81UjxgI65mUiOYW6ZMSCmVaNECliQ+Bba8Dgmm
clJTrbcelgsIISvBQEyku7TV3fzNlJQq/id5pKLwN+eNtA9vcs+03S/Uzt0cd4+VGo3gmuykcTXX
hkxSWBQBebcH2to1fzwIdkLndnFI1XrWHTvg46L44/iYVBJFoRyOVK32PeSfUUi5qKO45cqbZj1W
X1S8yJdBEEY2nVTMunI4gEme8SPpjy2riDnni0AqQMgdU1kOPXrTLNttkZ3RJaCdUm7pF58GNRAt
NNP5gaobXTQOlVRNwBIal4BcPvqnnxTucBN03/3snAk8kGijggERKKHnml2OQhwZmjEuSHntlt2X
x8nz5NfMClAHzG+EFP9XXhaCbrClgbgqZMif1dMLgDkv2rEvtp1toK203BfwhX2O7tuQ9ihpQxBW
0IuOELDujtmWRrvY3Ac2je7eeRcbKXjkyWB4xMsLSSOHTQhx5IO9hJ53u1gJzC2G5ah5Ns6Upi/5
yOoeqMaWFLSIVoAMyIUPkreVhv+gU5p04GL+eORJQr6Rn50GVrswooe/fiQhakKQMLSVDGoJEm2P
43WGTY6dup9sDkUoUzWOOsX6pHv8Tjja+v/mR6eVdb7RAywRDWAG2HQKBnaOn9YwXiuUvQ3Q/yWF
ypeTlLlQsnVmiRBF/OBm62vCywxsEafGceFGgsb40Pm1pNVvGdAQIrM7GM1Jn3Y0SrjOyUmxug2U
5vaGq0Y6GehyJ0RfFoJg2PboMJh4L8ELVHHiXDUo1A0iUpAo2XYKU7+3SfiTAVArJcfBcumw+taQ
YKeZHudKyJ2lRmkm3zq3VyGJI2LC1R7ToX/nhcf+aid7OWV4flpDD7a3esQOhhK2qqBhbkJOhlvo
v0hkaG5kwpqMjIfNnh5W5FExqUfpheM/hijUOIMsWiOGWD7o96aotIGkOeC+MoMNQ0N/aXrPnQVu
nI3IhC/bxoxf9d9uwU7LGAmnwwyca7qWhOLQrkQJ0DH294sb8HXyiTUrZo26Z/FjYandLiPYNMxI
ht+TmdAMAX4JahA4A2njN9TPI7C1qmSkLTaqVqDkMCZmSyIYPiKN+9izpexjejcFEgXrlG7Qrnud
GgRlENDMc6I+YOCx1BnFRA1hqZzMzdDV+iicLa6pYIgqRoN40dRLbxVKspJC0/yqlJE1Y4xp9YiN
AfnfODDdqwwRi9zZrmrUvUZ0yZJqVwvzsMANVeKgYsUm8xcCe04zY67cAclLM08K++aNCHn7f8NB
BodhOIsbPM5UVn8YpW0CpzCgKnk6s2Ns30YaXSOdcyW4cp07Q1W/ax3nmX3IIDxppd/WPAno2J8m
LOxrjZ9MdGZ/xE4xF11QzWjhizT/dv2MtUm1Qa/v7Pnt+9RV3ort/+zhf3xY6uXNxiuotJJt2FdY
TM6yc33g7iuBE9EhwITkZbbfkWkp+Ox5uAu5boSGxOX+YTZS12ny+pq+1N666NBHyOtvrXdHwU7f
3AFzaZtCUt1r2cUumkPJxOD7BxYeqtyg7JsN57xu09Zi51l6en4QQouEfoULerHudZYwqQqzDmip
JGL+XW++vIdMxOU7xdREg8Ovx465zLiQVPjB6S4eC1RBQF6dlRvIKBSeHiGPvTN3fMkLbGBrJGGl
4tNTHofBsJJmkVU2sOxYbpy6Al+XCASmkhiXFevJCWMjCy8d9pzIa/g5aU5+tenlB0a8UeeuV6Vg
OIt0wbpp0hWtDlz1Nc0L0tuFa22a1xUEw23zk7ad/OFgZ1NwIMXqWjIoOIPW16gWUNmVYpPfTQ8X
l3WnV19eNYDztIG2SXrRPE2TjIgplKhxXHaZNxxvqY3iI4Ug0W9Y57fi8oSZr6Q1Y1rslINaXc+Y
MCCoNiy9QCHCIf+ov6++qN32auLJbTpiP3arBcFXcAAa94DLiNcyr81cbXew9YAfFab0tWR3U4Vi
Z16C3RxRbXGti5KykzsKxIbLtWtDD8S02KIxp7H0ixV3thCoQHogrQa7Y0Kp24Mx41lMXJAr8GEQ
zKYsvtpAnvc7CqnyPbAKbSZz89O1r6ijQSb9Rb09jKjVNbeJF3ssuc/5Edw1bQlV7771QJpMfj1D
MqcgmDPYH/fwqU0/bwxhRyJiECsYojMkJFp0x6pHJw58ANxfJcAUt019oOsaov/6SvUVm2Ib9rox
Gn8FWmlneZPVie/PZWuHVOb85l1a8GB0rzrBExWBwvYsXdUIQhys/CqJbr7J2FlnJXQJlcN/wGhw
R517cwv7Dw4qnxT6HtMauWMezGFvF69dDiFTHvRKOb1ifRHcD+yTv9wgYY3StwVVYgGOnKQ8wNuQ
WD+R/PUN1t+aPNbpsjIrhMZ51+zbXffqyEB+9Aaz3yHEN9zB4xJi17e1PFe/HIckv2PMW9GA+Gu4
6D+1se8Ab2EVDEWoK0SXKuU7WR+ofrmjYd5kJfiqseEjLvIVkBFTZITn+nJyb1dd7VktSzxxihx2
EvH7w/nPLTDB7Lph/g9qZQuY8JMmndTC9fUXcjwro/2NADcdrVesme1EOuaF99waOoHPu2Hszr/T
Efvk0lvowR7FX7VGcqVfYo2XIYlodzw3wM8vhJ0mpmZAC77054oN+WVWKDF8nGmx/ejZM9uqLoKg
8ustQGaG+HexnpjMNEFM22LposXiniG994XYELWGqlmNVb/zaQKBHuziprMFu56s1irG4Ma69deP
qCo9e73QLbDSV9RzLNW6X3GmGUldjT4ONLh6dCWjBeD7Dxtf0Jjt/HOSfQPb69R0AKSmqAOeyKQN
skX/EjqZiODT+s5M5wsrgWL8xZm0hUJdFmCfzLPmu7FYBS+lN0ZZI7rN0KoYY1D5AC1xrPzMmGn0
0KkeYZBILnIEG3t/OkqnbV3tyk2LvhIjOUVnaaEqaZI3FhgkB/L3a3CUrXXsVyeZ3LJwvUg6H155
UtclWxC13IuebxtPQkfrLFZgVFStifcRCp0uAX0enhwSpmRFRUrvezni1pixSRqK7GMZL7e8VwZU
6uP0yaTP9r/kyclWZTAQEcJVRSrwgfaTIJjiESPXmbA3+k2Wwh/je8RrI6gGuGteXgq4FhJHapyc
Em4uYqU9TMdPyX1LhTCgHeHhsoxHzeyxQrufEvshAMz6iC3EFHq3PkkoWb+79RaUTl3zgt0+gX65
ol40ra9p2PhTTihQov49nHu9azKTLXuDnmbcknadeqicBgQx8BqKAgdeRYCx4BxgNLcgEAcHHaoL
FVYhigE7/JkrGXJ82tUD5AVLeTATfSP1QDfkqWl26S06BFTRD600D3DSYuGIISo/52Br1hTLkcx/
AJOBVO1XAdN/2PulHilH/stb/6S7fWeOQdVkqFQiF3z/dE00f6D7bJpGSZwq/Kym/AggbDtP/87L
Gdf5s9cTYCTHF+76/2IrQehM9A+WJKUlFDtzdvmZH+0AvhDT+5pgGD7rq3AUcCtLE7DyqO0AjeyR
fUFy7AbZd8gpD7LXg+oyBDpjUXqaXw7dmJyhWJCmdUQRhm2kSgKZ6ATHgm1Dt5xF3b4h+dhk5AxL
HXpv6BW/ACB+Iim/gnOHAe9DIkrU4Inp4gChx+TLaCXr2T3MVhhGDWj3B8/1eIzxZQcgnNmuvi3T
mokcCzcQqZI56iD0/e/B39ssLqYcBAswSjkKQ5dMmW6AFZKJe63GLzJy9vbrIjgTNP34n3GYMFfk
iuDPzJhaocgKlQeMRp0RRrdxWkLTIFl9SdLk58hN6Om94BTDAZpxjCCpi0TtW8A+DnA69YTAZikd
W/QY7M7SjuTxX4HO/IcqvmJuXjjM8rfEEFRRcESupGbjVCmknWGVKuu71l9c2dplyvG35SUQC/NB
5rf1KecE/5dPI9qiXlr2e94TwBRcB0cOA5UFShWi33COUlC6f3An/SA9LyV70bYUTynhoNlwpi0n
FLCWmk1hiqXqOY7GOJfnWiU4D0f/I9MVMxeZRHZzpQMJ+jjwl2DIn7iU85rWeJ46KFoREa8regG5
A5xtyaqmilEppRFlSX53wWmxrDJg49OfG9R7mbOf+zURwvvfXyaSmgZ+60TtjpdIpWPZ+WjUDitM
Lxw02kRfz9EnfveB0eil+Dc6YH+8xmx85Rmn/N+Pt+HtFUIa0RJNOghnxSztbm/RSh/MWkc/Uase
UqzR6uTwhM7a4Q5qmq+9I2ZFJSgPkH9vV1OD9XYUHcCiQ5tAoU1yGMPkvUvvraG6UZM8nw0KlxRb
B+VpdX39Djhm9hYHODeHNwxTvrldSCSgZw76GvgZPtDpie7ytgaVYtwo3JU/zhwZS992hqxXQvo8
Ne6VltJdOsz6k682kQBz1r+BPyYwFVFT3LdiXIanmhlhDQZuhtcmHzqgo08OGhMpF6biJlP+bJ7Z
qgoMeVfa3NFFRwN1mgOdpgAFF0y0b0xIjO5Q52tfJ0WfHaHqlr9cQnV15QTPWW9i+wKn/9Jd1i0G
UEjmyXAOUxjjWJZB/hl02dpkvswTvLb2ICcl8rlPpkgHbvYI2jZUaq7BpPqf5f4rYaXgbTknrtE7
OSLkeu4Uff5UK6rrajncd6cVyfkbLzQR8FnUHzapmSbzvgmG808MvAe5EwdRDtwXhx5fdrgfRS4d
l5fGXGGSDuqcX7HcRK1SkRYBwbgFKSMU8zYkQ5pXJLZ4gNB8vVOFIrfpfj36SM+Ir6eMgkcHMjRF
T2yIljIZzm2Osv/V68dgsoR68ZzymzaMzbOL7N2aYF/aPlb9OIJpBQr5F//JyE7jY8xpGbBeHvIU
7OdXdYwbeNHCvLlWGLKVNA569gXC3p7esJwGFh5Kd6GJ95dqwBle4hBvny6x5xJApFpY2lYgZIwO
IYLxywEBub/DwEoVhoX4J6gUnkbvhTFozS3XutD/+sTkkM+D+sPEtd/9+IqtM9jBevAAIHrP1ood
Eq+RmIXq4zgJbPJrUQvjwp2f0jwqIi7Hk1FpQl0E5adnGH6lX4qRPOB3hxm15cBbi8Uhy0oPLLwu
XvFvHsaFGIvbG8sNK5C2vuYkO+GTkv76LsiRA8ULUEH9Z6R5AiIX3ZgqY6APD2nb1VWcBCfxprls
9jY2fztzuLKOT1ZR0cjwKMGoXutKOTBC6rKLwvt7VDVM9h+eYYCHqPDZeJ5YL6aOHA7jUkze52Sc
CbN61xbUtcNf13HAWvVlSoSZcKRM+6kFNr83Ae2HniGkNM2hS0YkfQbxun5cSpNxKHsNAoiMM9T5
2eA+3DXr/bdDnnjP2HIkZpLtHU4KKOLsB2ZkumDZYu6/l6lT69TzU+Z6fPNbVBLP0tvrzzdu0mXH
4oU1UGdA2In1jEsANLbR/eii7OYGLvPJLfqywdIvC52fXMfD1DaOMHGc3ClISlgdHPzIv5zbWPKC
5JSlonYiu+V597DWta+yQaAjPWykdpnherzv0HYEWBNZeoC6FlRShH/Dsj0wAhaFt8+MCcAzEaXY
Pz+8YqUjThnx9hAiSdj4oE+bWjBKVDx2rEu5BjVmMc5WYSR2hRcYv6dhFuiW61V1oGfovBXAaW3L
yoA8PH0q0vSGFpEDDHcCPV9g1XKNbrdyJIW78MU2hW64QORkqrAj1smWmaj5ikYGN62Q8YGmbBBR
GfH63hD4OAulcDralq8vo6G6sYsqOt7Qzv1Vq5BHBRzzilkMISiktfhjr5WfR3pSgbBE3bEf/eWb
+777VwKdPo987YBeuT0HDRpXsexSr6uBithfcGE67Z77Ryd7XKSNFj/PbBmUPaaeA+ud9dw8PPvv
xa/blkXQkdR5OBxLU/1/oSfZtiQszHDlySPKF+MeLhH5R8heLlYnWO6HaVdLHFBveMgale1Te3ht
MtVAoMjHD0gitPJsJUrmFze0WbebifK9+nj4MASPcq8AVFxVKwwMkKvFdyP/MBaLj627nToTi0Xw
cMTScG9Qjs5+4i9UocUtNWnb0e1+oKz2QxLVGJBBUPnbnCOdkGP/hum0Dry6PQCakWxSFDiBggtg
hNzssZNok4GHly45iDN/NMoBZOCRjr7ICNTMTUQy+Pj8+f3lMp6cbLGZUzImw5iNKDONGfmPKNT8
CUHN7vRZIBrhO9riEU24fb+rO+spnqorNeQuAKG5Z7TpeHgxL6RT19JNPVNqVNDBYPYTUOfjpGX6
erL9l6mYBuJJB4tIAlYCOSuJy3EQqLoCU0q1Y2+vu57SYXyoJwSN/ZpJ2JOFgjFr8gLmL4RdpIzu
jevBlZZP1Yi7UaW63IGFuQVm9e/+EeO91J0/iuYCjWQ/1JWYPdDUyx0ttnVPp1Ra/QsPzvG5qQ8c
K0+sHlSv2VRNd3srAGPJUjTr7sNJOantEEJmOTQKtjnGtBHw/Olzk1KiqwuEemGnFnYCBLXed3lZ
5U60B2irEelX0aiAmXLYr1bpkFR8kloGudtAdBSwHlfHqRtLcSW7GORNslt2B4wuT0Oj97tT4msv
tNgg4OTwChz5k7RILF83B9DqplNDUMoZxzJ3ZwksAl2jCB1eHDCal92PMvlmI9gAxNdqN68Ea3HE
YUPhzAAwRydpo09lBlybsSdKfuHppp6hFEq0sR+Kj2/RBr6m0T5kpokRC3zo8Gt5Cbq34YfexhiS
NcwkOIGXGCYsD7mumKQ6Rm5tk/M+jhTYhh3iVIdwwonGZsStj77ZCdxBF57M248upunS2R2XWAgw
hen4gEew2U8YwevqUBjBIoKAmZRayjNJLB76L/czLRVxYhDy5F0YZrle5X39/ltfC0NP5okqu11Q
jUI/7i/76ZPjOtF8JYY8sjQwbO+/SAoESBEbeMbZ5gmul8c9gyggi5yKSna92rUBntjTWw3hvTyK
3VQdF37NRlcLd5Yez0dzN9cxnDjnVhk72kqxSPcRIFDJtH3szZFf3XEK2zoyVzNdYM+do2g0JSCN
dG94PH0kdVmKdmIPmkriBFBqZ6mHNPCYfF/CJbeT9fKxdm/XSLYhtLeStCW9gjzD6HRpVWECq2js
iQhsweORYQYgqdog8A5oV6ZOogKCHsT0pfJfpCaW9feHPYr0HM/6aXu3FTREZOFsYEp2cNf7VhBk
Lmp86dK9FO0On1zGF6bwrjw+ZuFR/dpY+I+si9GIivPOmrH8VKhzEpkZgV0A16Ohnk873xA5C+Z6
sHNTfqd3Mxsiin9us5qIopZfwaeunEbBqiCDHF4L3cPqVEpA0HASWy17OF6xV3aFmx0dDWDMlPzP
MPYVQFILtp6XPfbdIQgEJUCtMDxro1QlMERBEgbw+BN1Nmy979yUUZKX3FydXdu+XbL6ucyRuz8c
ZvUNDcwg0JP5inNJddJt3tLJx5AzwXIfwkW37LOgKvEMKbzMT++vdawYeX+Aj2Id4tOHNFWtIKCs
K/jjQjNFgAtV5T7eekalSol8HRyVc7k59q03nROUu9d5APalZdtKPJGZN9ErKgdD0/WuVyePvtMc
gxjs4NaObcZOyHAlFvya7b0swlYD0V0oPN0QgykYc85TMB7GgQYl017fXXyJPV3gNY3QUQpiibGh
0W5T02AFo7pXckPcMUCCFPx5KKd8CmlJvSl0CycfVqpTZfkRQe8xpgjepUNRB5hrHxFe0LBG/Q9Q
Tq4xwkUM+i3luZ4PYz9J7tcuZnUB5HRnpWFfOTSzs46/eL/6v8Y3jSwFtwW4Zd/AXmGFkGOXYWHf
SBYWjaLffrEBymghXuzdUK9CIvfCCHUmv7VANxEwDQmkRa8V51zbr4IbnTOQ2zjSo3InYdG/rGCl
mcBTo3O02fcPSHc35NvzIrwIKukrNaLN37d0MeokyeY6Ttt+FbZixktHYm2ta4O0m4xcB51AD+cM
4nMsnm5gA0bBeuhimUQEob9ciG+PFdxSriG69UH7dXecFs36wVtcVfGTcdsP2v58C7xOR4qcBu1W
EIlB6ngc84o9zIg74FcsPCxkvlEbggipd1dgBLuqGiGLjeZDekfsyxJoH97UVPZya1DIqnlixIjA
+CIiqnQFypzksdz3YMPAh0UmiFo0fac4CFbeQZS3ffNUagSW+SkLNaZuPP6uk4LBKVa10AXlVN+A
z+HW0hPa1WHUhi/zKPZmdKO+K9jxgvB019QcXtgZEq2Aq/rHqdfNTh8Q/wW4vV0sBt7m8j921/0R
DbYnK8wdzMhdGvwHsI3bwqiPDet6/e5EwS7Ym9LtR88MOBVIqcIB1XbL+LYyGrkpIhb6C6Ha3s4c
EnW9+Ia+88/vS74qMBL+y1t5djvUs+Q/K8RM3/glv/Iq8bKkBcnjSwvtEiX8DkR/iLcYhxSp/5l2
YkGGPb5w2cEtmRa8Im8mAG5U/hwI1EiSJp0MXSPQR+fWHXRDqh5vy+uwrAEzDsluNTLtvCDJOAco
VM7GkuI6E7MwOywBaPshQKX36P/zvuqm+705Z4yRnZmevM28n5TE/PO+mk7o24YDxNi+plwTzQkj
ErLLCnl6rCRDsT+ZzNqCSdGTfcbPEkRYhz/FhFtVS2zP/bi1oaHdp6LA9R5RCwvvbCLacprD7J3/
gzF6836e05bEj1bnpz5itFjHSLYwjepNBDd4LofemEuzBfPI3LmtmXf7wxRWOp3TsP1g5gqk+6vU
yIUlhrTNrhCoLMKAuBxIET7BcNiJxy8VKTsjumrb3lNvDLwXEp7dU6Fa6SlZOV0ciWMnyJ9KtDR1
JWf6nkhurgyCWpA45VboAzl8SBupfhqVGCEK5Scmz9JNN/ntWfzOgsW8ib8H3zwtX45lIxiSeNAi
Ee2Hdx+BlP7Onj5Q5BbTDK6BmzhjGrWbTp+ID+BewzLQAnAmSzphpj0QKX47ESrULjEb3xAjxIgZ
zadOloMr+75kYD0xliwP9D+Zqpa/dgVJ5HXH9+JREsmO97Ns954nuXfqjEMXTvPgKqa9oOeEPBRX
2zQmGppZ7aaRmbPMumBWqLscsqrB0MvEHGN3AUvGKBmFfpgyuD6c2eqjzoZQtjj2WCeZ7LvazITq
lKOOLw/6IiteNi/HTXc/d/wYbXYJ1pXMmo8MPgmNLu/hP8AoCZAlUPeCuijrKkrM5IhnHZai7AuS
gDdcAXhQtJbW1jApDl94Jknd/rzBK3Mp+YttfjEOWyCtAxsB2HQhdmcGZ6E4vegziCIYW9Te2Fug
bS59CThAAxc5sScc0Kyed/MXjv4Q8bQ/u9GV7mV3gR1ilK6LTETnbWUprYnlRnGM/LCJ8UZi/r7d
xod4tioW9BJStnegDu6nfyS2iKD8vDD6dLC1UjyoRSeqQ9F4Y1ezWB6fnWta6BVNGoCOTTwFG/Rg
9rHPw8xndxNTRxRpU79GEUHCNd1dNpzFl0NnjcaPHF52SD+qlUeuXQbE+W5L3rHe2rax+N/+E1u7
g2mj1GpJud70z9UN9VD76iDsWj74NyB/gsdOjRJpBg+Aw2j+Vj4v1/aefyu7c9TbOAxtCY75RLgt
Fw3BOi3YriXbrZZJUWuQyhnJGWCvCK1ahRYU1/vLZpHRS2GOPEWfIR/hru6EZQ5Mhr0a2tjxGMSo
qT/UxIxNm/T2lSVXeUYk9bR7quSJqnuvv/PJxdIknS2VGX7rvWdGTWhblWX7XtYawA6JmCjAaAq0
2I3J020kWfgQ4eok0egF4pEtqahF16QHR2JTqPdMN6ty4NS14kkNXOYJ+VXbJuokLH90QNNAdBSY
8OevUmzcJS7ys/IkMhKKcjWYy6Ndbnb2YxbILHTzy7C3Rp0DNjKS3o5Wws44DRUzsbrAmTkczmvC
BN0ayb3tp5GncF/HwgqH2Uz1AbBP48efoqo1wjTLmV9oN9klHCyGL/aBL1dtgIzI57Zntt7ei7KE
r0IxvevBLlr9BMr3A0fBdImHdrj5/kSprvE03TIQRtopJtjVVVHjcutznGc5Nq69yIMXZxh2d7Va
Wb9eRmsYQbk97z5SrBbqWsPbHzdIVBtDSeeAh2is/7AJqyht0psWsmh7klS3YiLetP6QZceQx4Vu
3h3KBZdI1zPvu3vvGVqq0JRE4qKXjy6JMrUfVDWNe0zfdx04BwMnKE5MOlNzKaSYNGS143/lrQ9s
R+6LzTpVozdSaoIYSwHfOFT+3GuOJQNze0586BtpzEYqTlawUu5EfH17D+golKjxSwG72T+CYGEL
OSnJCnjOpKXPU5Zc/MscQYmMMBta3FhNISIp2G7O7ujdZLfJCjFF4IEo7NEkMfu2xtiMSqdBtS5u
HsT15eIkvCawCff2L9yROSqe7Uu8sPlKHKbofKkpd46Flah1rAoitHOCPLzPeDmRXo6ocY0WtWPf
gqktanaxjAimz6RU/dMtfdIqZHcT2Kjp9EEGtfjbXiVZ/nTiKpAFQuBc1ygbw2n9AuSCXgfDNije
r0ym5NTikc20+a5b9IVNRFE/f6yhVm5YSEp3rIqT9YBsXv6mlxbYS3C3gWzwFevPwMncdIKpZ4UA
S42Hvwa3EkKV0cwimJzLoFtXIhwSgFhsyDg/ET/GjapWeFT4brePev8jkjvt13447h/Wxu1INqxM
zVH+PZtJMTUDnG48R4h23jtLR0Ra9C5v/6JyIA6PWAC3gbwkUSu57gc3cWo0YHGLzpVEuIBWSq2o
3N+c8KvJTDu2/FXBEGMGaHaCgI2gpgBcQyIr2hitK0RGMx0Lz/BpN9Flk5Bjuop1jUzU/+7DlKUi
zuRCl07nkMQK0DkMmoWbZExTqrL8UrGq2pAuE27Ew/H58gL1iThWPCHZbUDFXAOYwTJR8uloMFBx
Ivv54DgWTHqPyCrnzqV+taymFvT4mb219CC3yzs8boUGCMv51oDO3OE37idy2QLnHjE9Te8pF+hq
sVVLCYTu7j9geibjQ7oEsgfVWsVVguAY8sGjoGRLeSZrxuOdINqdWzjTgdU8cc4gdsGkgS6pI8VC
+EXhCqtneP8N0SHUoRepStG11LXvSYYj4R2eLYSgO9gKbdZGE/9TRDzKFXeWgkjZp7lWl4YJmZy+
71KlF2s/9qT6mtQZgO6NvjaR64yq7IMtv5xtThhNoSg0D3p0160ANJpDQ1ZSg8SxVf0BOe/LhRa4
34wdAMouEvYy6/kr7o3fhTSgEf9mp77rS9M10TRRqQgzOVMNhT/3cglYTPvwkdIMFjzOy2wYBIig
uZOTTKa08+HBdpo6JJ7CDL9M58ivy39vFCxXTTXedY39H7mi6ttIUKnYEqNi4VNmnc2qVg86sChI
eDd3mm/o9TexuXuZob7w0ZtTNuJ7H2IuecUrpFMM7VdVMBF3FhYL9e6J4t0WtVO+MWSKlHfv+wnV
SjueKsLCCzNpEjiPf4nog8sUNF360FZuIUYRy5Mm5Cc5ILpAdx9GirXD8bjfxq1wwY7dcLq7CRLC
XbXlEKy6cksmAG8tFbRiJ93V+KW3eGOx7dwi6kA3R6t2+0TabAHi8HovydxpFEnm9TmGsJjfXAnX
Z1ZP42OclzJG42Megle4aeeptvnuif/cc97lHwFYox3SaJYVj+39Dw8upnxbYWsJRiN0vD9MYzI5
ZmwdUrQ6mbkadnuagPKCy5I8WXrDKEfm43lceRWgoiMNiBZ7Ywy/O5PUDBw7kB6ZPd+/PUdVRLTt
XuTYt4tFgKfRkW4eDGT0wFUD5FeKKnVK2GC4MWmrIBuwve9WAXK9urWRqMcuh/hPKrIFUPpByqeR
9Tpkbc9jaW7yKbgx1lrCCkXKzPN99xqj+wzzeBDE5NFZxriZ4v01gAv4oM1g1yxd1jpuV4NYwWmi
dava4nS1T5yLy22aOXCaS7eEDI6xEkmE6hT+pgTefpl++3NVCTmgtb1C1LP/aef4dkofo9LvCI9A
qjF6WqA2FEkmMI5byyRAeajPQWYDj55Iv0w4/ksDYmeEnE0ICssK9ss7ZONWGvYFhp70/GMJshMK
byFfssLFRmjq6kpYdIWsvitnHce56mpMfY33Z6zcgaam1pSaBpWiMNUo0AG6bTYuoHuC3MHFzfUR
OaJBRCM0LzT48aRPmf2bRFvFd0VPE0LiuAAIpn/8M/2TG62daLCiOyFgYw9kQrfBPg0swkNS+QNY
VsKGlhq8SASQKAGK3v1uBr95R/JrFCrO67fWI0u5MQqPHNgHLSlTMnttUKAuMKbe9ArJ6dof5yiV
KmEWR4KtOE0R9Mju6wsKU6+nAhrfTBNAGepcyMQM35ohbFkBKj4dhCQp+MdH7b3n/sanO7SWCebf
Xqid+xmfScZk4XnniVBmOYSFVY+8uAjUKn+gUaFOAea/vE0KptWhGpX5IPTAFaOTvgqb8Nb/e4zT
g1trg6IthEYYNLnrCjbyi1WOxWA+MqbsIXTiNIhW3Hs5pjyOajT8KnjYxZ4dRhL1vKPo1zCYx+Zk
y+PAdIRUHD3tLTIhLiImRRZYnVYiO8elQ1uIYzeOHGW9CZSFvIZrX7qZYK9IIrZSehyJclXK22gi
rEcVEBchVXA4V8C53ZbVZT9K+YCRWZcuAg31KSv8hhoBq03zT8HZGtuyWcwA71Vtwc5+HeXwtnMj
27TvbNpK0ReZ7zUB6kr6idp8L8h8ttIo5H8j3a+mOPiSdFRhopbLmDWRzPa4tMyJle/AHYU5cOLI
cDS2swo8EoFcAbYAlABmZJVBsJD6Vt5OpVk4ISK/UOLSPAhT96ooi83aKrlQAWWvw38kNAE+T1Gx
Ia5heImdC3rApWkZhExK/f9YSiz+62FMFzeYCxpxAboWBNzR82cMdlZScdjg+1JHtDxqVzZS9Qci
Mp317p5J27PsdGPBlxmO09Jxtqah+1JKrwEEjMAsT0Q3mxqeJHHPisNtixuH3jbFxt4xko1Z9C2c
4OMQkPY+0C98pRPiS3TFpyLkVJlQuHbMdTu2D2+iC3cCLbNAKdrb9oG7JVeL73w5ppBjNW0De40X
xl7WdG7qEU6bPcCztTiEMdQVMm0RqFdGyRUih+fzKQ73+oR9oQeBoUaptDpw13nvVtNuleRj57Pg
SDDs9HSvCEFl32chhEFDGCF/+v6w6Ie+2JvaQENbI+hIT2LtpPB1/8QhTC0c+cjiZoyGhM4/L+Rj
tN276t0wR0x9EC97vjnHlLHjccL+5h4iIiA+hLXP52F+F44KWRnvZwD4ZO7IMsDIkb1nsu3B1zF2
8KG/SJPGZLW+T9XwO7JkdH5XnPH25JQG2ftVSkvyga7O+yIoL/Cg0RKXSsGYE3R1v8JRTeOhZ215
YnveMYD8boXL4QVNEB1dgPDH0AVf+IQoxxBRoHo4mPi8GqH742KVhauQOY4xuoQZv758A+UJDhgd
7izStYWRNlXX5x1pePtU4I2MD+gbhi2nyNJboN+yuy8bMU02/i0eyz9izR5P6p8rmdY7YUAsJT+K
RpYlADUh7L/9+UB67W+FU2m7mUm2DNM7/8v7sJh8NHxt9amFuqoe/iN2tK1eUwQdOC8iZhL/pMyu
RcLf0ywW4DSrZNFRnbi96WemwCpNvjXubUrBsJ4fwfXMB7d+EOWkgxJ2nYFy5XgjRnOgAJWOIhPB
owCTJnmtnP8hgU/hygAV4DrHtEBW0VgNhsidJYwoSX0epEVBhvRHHsIJBqKb83wwyoCjOOUrkswE
+zHS/77EKA7szMoux7mQvtD2lRsajci3RJZx0dWMorZHu//i1bcpKeCQnze1sglIZix8B2DPgYDC
QxODh6XFChHTmmrbrZltbZwwkfIfVu4OfycYeTxUCtdD7OcGLRfjgPdnO47GAE3bh5ol0KyEL8rn
7OZeD5jYeo0mzHQiwdlgpBQA7nIB4GWP54B47r3pQTQ13MqHIG61UnyLcN68Se7yatr+0PkAjL5U
QaJsi2ZbOiq5K5Xt+CbcGObYWf8ZpkKaFWh+XnNAcxk1rUYt62KrO1RdgcRNfIZupWN7nBJf+SzT
IOQvZFAGAyXEkuke9Fq/ke1qNREY1GGpUCBHDcqrTgDtTyTTNP6EIuLyQ7q08z04ERod2Z/jXsOj
audoY9w4lToySrnF6V9N9Yd+4+/54TUmkAvvR2zOp7zz2DF61gEXOr9J6VgEgGblLQHFrwYTvImz
mg8BOwMQO3DgrQvzGua0x7Y3sWvWoMcPVzUU0Fo/90mLaQscqXmgjuNbWJDP3CG68h/yfurZY0QG
PUlVLrrkf/d1jNzdC1OMsDXBpSfDQCIfAOwiwiYNLEKS7s8a65BwumD/RtT0ljw6ZQ46Go3cNwcL
WdN5KzeFIMKxl5OBMLiIU0Hh4shPm/1B+94ry7Dd9GbazDlisw+ZE1BOfwjyehOYDG4jJ/BJOGpR
SCyKt5rk2xqecX92yFRRbm39xPqYd6OO8xKU4VhqTW5cJ905l5FOuxT3+/tnNlzJS9KOmf07GgwX
OV23UibxdLIRBcTTd4ZUo1RnQNGr+483ibYMcp/R87iNYyHVu3fWRBnEGdCfUP1/dXlzit0oZeTx
AthbFZH9mHdklrcnWmwNeiwKEFxTmgry9c4bxHZgmnbno3yjf2yU93BD4KcAm2HuIdmBzZdKFO0l
equtgbcM3ryttetS7K/JtgagPKbFLzp97gF3s2pgByW38p23zaA0D6uoAfGw2wBzt//EzxpJMsfA
TkfS8amB3m1QvKKqfRIxB66gA6vJQ4WOKisiTPH50ZC8tQZq/nQ+2Dfc5NglqRo8FLbQwnqE0VZi
zPW5YrOpTizwUuos1amR3SSHpLNlrXxEzPRUn9DmrJLT7kj3AH6Udt8pK3zVunkJTqdxLkdsJA0j
d77qxJrmYkz+PG8YpuRIMbSPGuQKwYtkrV1biYI5stYQ9TMsAhiWH22Bz4XKElyVBhTSw4oFLpbn
Z98ppmOF1GiVKS7Fz7iztT7njSR2t/azMPsBm2XqVlmJfHjb/C8dxfjP4+MgDJlGhG0J2V7n0opH
xMWLmkEl9SDuLiRZ0FmlsReaSKuuSjh8RRUbB7Lyn3ntgPDAUjCImYmud2H1Xmc19Jm3/knHD16u
diJtr2RPBZDMXI73y4BJLPbY8mhE7ktGmQe+wscasH5QtmVmA4Db26BZ9aw2hO9dZHyhYeIeh/x/
FBnBOc7BKcWlbW53lWa2Pmt+nO36e3l/dL/u7+PE0v/5ge4nid94YB3kf1wBOoAgIiFFMUF3X1U8
k4sJmDcScLImy7fCwBeQi0bEhZE07tDxBmfVM+xmHTnomV3mb94b2BvD0SiLnBGrJ5fqKRNCqx7y
M7r1ViixDc/xKq34SYUHa8wxhXhxrXb2Kt2zmr7ToEO7giPg8VXtrydSriR1cgcA2T8TkrMbl+K4
7R/l+RJheBxeOX46MJv5s+ON+JOCVeE23y7E8+wUY9mvAaNlkj/fhNnxFJMvZRq4QvKcsg5se4c0
dkIu4phGE4ebBzkOssOJW3sVoRaIKizAyDSLw8AphpeW3g8/I5wvj+//IYMZDzKvYcnwlLc4sSe5
FPumnkM+aeBJ/I3iSG5q2IFy77BceG1l1W8qEG71XkPWU8Ud4QpMg4v/phZxFBn+nQIJTlmIBn8H
Oc/ebai13AoasQ/x5O4OuZI3mD5EiZ7H+HnRJRFEWPK8FEegX95aGlA38MMG/QWq8rWlObvcNjmg
U2GDP8ae5AEyc2cMn3B4cdFnSCrjNhih/Y9802F29pRbw06agkYGzRy2wBA+ZG/YpgKDGLK9EJa+
dhh1fIqzTiiBjZbBA6c4VRlYecGc/zlcm5K4zHf+nyaMZJk1ICFo1Wc1KwublJ6vJ9kBbI0RzN9g
INdVwWFjxgduY7bqW+cZMaOz8OlwWGNwTt+K+RJeO9yIE5t+1d+J6qO3iCEc+aXkBbphlfbbstnr
s6kp22opJ50k3g1zNYBuMEWFwz39YSJO6KEOPx/0Kbha0PWeFHBAIYUdwriA/BcnzBZsXXd5dIX2
0nYshdST+wupW01SXnajzoKRZVHudNz5BiP77jdT2HrCZayEOmXCu9sQnHhpZmgvfHNbM2XgumF6
T1S4OesieE95jp2RYAoSp4hJZVSxDsHvGeovnX4tHx47EuBlgTVkVy4o7XKCZ9jd+hMkvKdBVBa1
An3dF+wSZaKlmx4vXd6luYY6D0Ox+SfGILEIZeUJWic08MrxEzfCc7Bwj6rkRgNHyytlhOqtmsJO
mN6q/37qfBdF3KyngHZoDPtVXuT4URJjB6+oA+xyhvExm6S0ckxW2Fgj1Z4dkuwEAsRPJIv/3q5N
wUjAoZGckL9EXBv469EdpNn6uWKeWY1yh5VMmmr8friJnAHEeMtGh++6d1IjWbjcs/2LzHkJizo7
9Mksh4AnqLkV6t6CNcIPbKwjHx+1T5ekmPyr5ziSzN6627NuqyNfx2s/VpD3Bblw5gIvaM0VzTL8
wOBEUk2jKYakOwtyEJZE6RZQlTui7lUrQ+olqaq6+7wWshEiM1lFyfmqX1/XXyOygky+KYom86/E
kLGD9oCxne25/t5AiGVpcw1IlKNcv+CMZ7+2kYrt1SJJhg5RJ97RUr3ogda2s+BXvI/dwLYPT/4Q
v+1w36n1OnmjeHFi2ICNGtbQ9wlZa313BiVZwOIRRktwCwrLAHt9eW3v/L+xZ63ScDA7eGzriM7c
82pL1Lh9vSEt+DZwiAJSp9WVkNbdp3xtTBR9K+h6xm7D99YIqVdGnShG1hZT7t4Aol/zNDOJrQYA
snMFtlBA/cvSq9+bx8KtBLMjAOZLBdZaPbKiMllQ4rPy+nJkvO2sDqAK8iNEMSapku3cgSRM1fVp
dNqdAaOttK3rCF+gtnNI2T4GdfK7F0XNohr3rldaGvRkmdY97eJPvn4lf/51+vQwXElsBbIY0RME
+7vz2JL0Dvrb7P9uclI21Wdt+U2MLxEgeucA7iwSbR5eT1RXYa/5BxCH141+LW4dadiixC746fS1
IrvuEfwyFHb7TmSihRs5yD3HnLz5mND20OKW59XySO5qVQCP1fy+IpIeveUlsaN0Xz0MwHMlSx6Y
5xmEHfcs3Ja+WgCb6+y7q3+L4prmwfZfPD0jzS2zGHDDH9XOLOYJJzjbJ+m7+mOV2kR2AZ6Oi8r1
0pE3xQbGAJv3O4Jcg01RVeKTMyIaGzadVtkyqdJjCoEfPzy3i8xgQf7zxFMrdzVKomB7eEYagnya
GSujP45dCXrNorbBOPpiP/2sSUQeuyXPSwp+DrnSeGZ4S7RUJhksOI0QWmyuxnqlHlxvfGg0ML0+
T12su9DTpl6VqgtQk1fiYVLm+vuOPSBhvOp5xMlfwGIHuU4FCJYikRSsVkXcvIMwud6PH38ggTm5
suwUQDT/T9QldcO5LGw2QZAYjlVh33vwEy4cAGSfkSCEkNIbQJWzAo7LWESryfav4veOC/WsNhR8
/0ENTMdELBJsKTJyosg0WZVnjQseYuifcNiZhNTH9LM6a/moEhidZszqqsFrN+DsGxctrVZA1oNj
NXpazTcCbhBlU8N9zOPHCYjZLPLFaBd2ZPTuACV3hj7KhzQdUymdnXAkRq3VSJ5cdosYC4ZLIPZ8
PiicdlS8OXBN0a05pWZF3S15RnvLyg1eRHNJiykIPIQCzZVvjC5BmsZcL6dXddiVcXUMSAe1lj3e
1iXBGie/kOLpJgNDbfhgn6Nm8NTAIDniiT0osiEepcCLMW6ZvBMHi+Ujau3Iz6qZ9+KqRFRAQ+++
GU8KPR7tNBdY9Mc6sLOn1H6182S+h5VZbGiu+yzh3pvy/h+YMFnBz02YQ0A7YjeI6rWKgRALRsh3
lFL4QGLLcFo3RPom7+9i5CaW753zTt5mQnhX2UkfFv2u7PXpRElBAl3//R3GeEIN3TPN9x6kTsHF
OeRfvhhT/L5NjMRuZqv0gcIOgi7QwICAgr3n9nTHCgSqnqO7i7eDkCCciq2LhEc3pQ5RfTlIjsfx
083TTAHF9MstBXPDli8jWr+0Zlx3TZDtpndl3mkTwxIhBLS7v0gRKArW0vOWh/N4khjXOnnsDlUI
WPPYD3YHmpmswCbIPX9usoT7Rv6o5TPTQ9TyNHRnnRTcoXy5SV6PXxZPGD0ucxqEZ9jlCrGGxqEk
NXTtik0h+EueRWnLxGQ43ZWelncxGwVOsYJfbrQWugmzeLnSLMYyYVOvz+ESOhd9Mz6M19hXf/ys
RE/RsS5kNH9AZsA8VQH/xxfeGGNtEmuIgoSmHaWoQnhwFHMQ4HNxvaeYT0p7QCztXviRtmpxgatD
uGZP99UR1qNK5tYnSMy9JA7r2+I1G9D8KH2KJbvS5cJRYGRmBa5RRaIOr/wn+utQiDoetd32KPLt
Uc9UKbNDBtISL8D2oum9JjLXLUJiytTq28GH3A38MG4zbjJVnm9wvP7/rXiy7obtUjoURjk2vlG9
vYpas1J7iNg5J5/5VI9n+ev06aseFTM57iH3p4lesmNG/CY1jQTm4n/CLhkq+kB67/NFT1B5K1Bh
cXtJcCs6LWuLheYe181UQsuUk7sKeMpsrMW23yq7qM3ET4xZPkh8N0NG1u7sjUMQNVpZn3og5WM2
qXdl5HeRcCMVEPpjfHbJaaIG32/DihEPcofCwsE2KZTRoUP7mj1mcIVy7oO46Lg1oxe7WIJbpJhP
paOso/pL5RuoVsP5hiIyZV/HrxsMpnedpgy+E+7V5t+AHsQUwrkib96oTHIgUXk2COqS4FeNbI+m
vHzl5wp1KG/R6kjXU4Ox/gWwHr9cDRYB0IrETpGaqi0kSxzoXFpirn3ShDu2SQ6mG5WYzQ8bbTaU
SY0cdIptmKqEYNp2jMeHvXueG5U94aPxxeqsw+6jvONa/8K1VnjxtM2kn4DM7mCmje9vvJZsGXhA
2cR6OJUpxdomk3ij2Co5M3j1etWza+XxQ8P3RAqvgoMWc/2c4EkCG/gW6sIjNRrOrOQ28X7GDkbN
S2dHHTInOtScX9Fk1sx/ptR9KX/BLJaDqKxzx5M0gx6rUi9/5xJHQpu48lfUh7UJOn0uTSE4yZKY
CHos21NH7P9wwZsmWVzsxXUGHnBdFjWntdcfet/7T1Uz0WWxvv9RTz8TrAqenKyhz8S9yQaUDSHq
tFG3AECakhDV5kTPZjkEefS/vv9IFIGvTInWWDc5l4zXTlGveK5S+Nz7O3Tic1QUFxs2yyynG//u
i6K1NMUdbrv/Ao5K2X72avXKPnQh1XqoK/nSzbQ7NWkWUsPPWB15/W8af4YihUeIQ/wXnkyEDpMR
TIPdYNl6Q/QZ24Db2obT/2B7lbybzrN4A94jFtqxHPr5rlRZ+MWkMmdUB1FxNu9uywbbtUt/kQ78
o9/0Yy8gpSzXxynzPMqLWnm2YBZWWRoKMxsi30bm+KFFBSvNJ2Bjr8kX/MjVUKkZTa4yalGsWos/
dbx116yteCb4oBKLhyXwCAZFpOIXVxyLDQKt9dmL7kmpb85zgAaAnLrk6aDaAaJIRvleBu2k7KZz
5Vpq3SJ2cRWr9YmUJlQdlE5MNQkinFnOmEWXwoT7XvFCDibbkUuDeqIUtf+TIQcEF9RnzlczksYl
Jg9AuLwLYUhClmFkwAK1XHNNuH9R7jbI9UtG2SAGo1FNwEopjJkWmH8CwCYWYqvQxgrMjTdzKV8+
rYAuKdXg4AcLFlYIGdRWcB2CAkmuutIA70LMVmyieSHqDpHR/7pj/b52DZYB7XQHpzMnJdHzFcdL
g8KQzyd0oBguDT8238qsvwucgk7+l9vzQdx95s30ZFw9OkP1PGjd5QoXIEiRT7UdON7S7bbB4vjH
tNdFTeqafr1UDpdMQD99iIqiiRKcGp37UsDh+cIkZ4++rH6FYOnY9yr6k/1lgIuQdiV+wIWpXs6G
3J1hUv+vwRoxd7ilYNTerpodlUZS1wPS6cob5P54oTgk4Utb0407KtSoFKHLtDCy1W5ZY/oubwDB
e166LsCrjqJcQLlLApvIzPjeyQVz9nMf8yH2dNEx7wWe3beYBaHWnfqyBqrCSXiZNBfqq4StWybn
5Ze3913KTYBX0gaYLU62Ms/60lsVHrVx2kcHlsFgjP9ASl9J1wAa+Jx7CfGb1QT1OcUCw+IwaKiH
tKQBJasJPIygjzy6XmNCOwjr2vs/fftxBFUZerH9O/6TjE3rvh3iIzE5zcMUx/tp+VWpDar+oN+j
ylAqZVvmyX6vgHpNS/OaKlYWdm1POxAfqJLEiiW82XLP5neXP+f42dDGQopwbB4ndfXmWZs7lPuj
F91s1SXe1jHz1Q1hqCWb5ktJ3ZkZzDqiZcPX7e3sIZRjPBev1rGto00lGfNvqty65eLVyJAnXpX+
yeZ6eUrdQBi3W8V1BeLchgVOFKPts4RRMIFTuEBvwlQENlgcPcNB5zjuU+z7vlzcZ+NRJS7Sp/rA
zHe4L4d7HtupK6tjEGEYwRmFvhy+WEviAXQd/1evPu1MBeS3a/uXKXg+nkc8pGTMkgIz+d2j3JnN
yPAa1B+GGAQ8GKX6dkw2rnahefOXsHId9Xot6HbI99bba9pBWsDDLXQ600J4/bfxiWz85jcwHp9m
LhZZ+05w27ojz9C1eSI+3FWceivOmOq8gibzC8JiOJGXW5XfU4eKylX8VIKn7JyLzP0AcGuHXo96
loUZXs/fUN7Gj6dIuoLYXWpIndCJ5UyIuddiiXIndlyEFyAB1I87jpmZdZenakQlF27FndxnN4tV
q6SVlmAoFgUZ6vXNThCPGrRl+clmPC2+3ToZuvQ14+Hkybj0oPCZYRGH4YT57CrpLZ2Mz3b5tMKE
C+Cj9TsGNjXoRezNeKRLvUJj7RfXPgm6AR7Ph30FyYCJ3kRX2RjXwyl3W9HqxN9Zmx9AJOSWcbKm
4aewrUtePkM2H6CNiGVY/jieLWzoCg+tY8AeGh+3qv3nvYVEc+uJNnYJ16xBrOIMa7uPgKYPWq9r
VupokuYVcnqXS1FrkQK12ovMtTynkcdbMUqHukJOCz0kR1Nqb8BQ4AfSE0UN5v+ZK02GtgOWDuNr
6AkmrgYpj3tCVUl50wHUvgKG624/uvw2JVh2vUuZgT/5v/Yjj8iehz8pi9Tb/R2ELHFPB8w9Wt2I
j864BUyyKSDeOocPxYVQ8gc/2A/CrneBqL3551d0RvoSElbcY/yZDplxUAkrP/S22NF61Qr/I+WH
HkGTfev+UbyMDzuE8Et85C/HDLegV6AhpKLFiN140OSBDRvUD7K4zXXxo2Cl/xj9ubqUY6/8fz4D
nU6KaUkwtsB2yy7nKLTHHKxcTGAzyEtG17spbJ40pnA6cWxnoqRAMSwAo9PVu1YwV4MW7g3Cvf63
e/q9YzwkXCXmrV1LNSLZ5jDjwQAWJgTa+xdvsuIPCD8dLSG7mQ/Sc1MejG8UzflYFUgptZqsO2Qq
sgAlKOBybBg8mzFd94VuHF39zv/ekMlduePCymvBkDwR9Ow1QKNn8cK1Q5uKR5AH58QdL39FxHU7
nzzl8lOkTps9THA1iik5ghS2rBAUuXsufFLk5bGa/bDstoCYPcaK0N2Z0chO7CCRbKZOIwzpD0Ub
14F6Y9ebmju2SjcMJDEDLBo/OaKj2MI/SWFbzE95rB+HgsdCaZpzew+fRU211KZTdxyDlmF2G6Ov
9Njq6nkJsO0ve+KafIJjiBmKBfAi7kJifBIkCLJSuIwQYq4HRWl5LLauV/utJ+FWChozpHQ17vre
J+SIRexzr84hjJU86Ku2C7lJ5XVTB2WwBzWmGgXMRUzWypLE0Mcg1hLOZwV0uOXYljC3mr6kixpp
LUVOK0DLxlFeQ6UQY9rK/rOWLQBIiSo9sN+ngXvPCazCLynXqiDzIm3UlnXB1Cpbvi9d5dPoixLq
lrcPW2Eu52GXaUkBK79+Tg+ePtjZEXOLXuNGOnMv6Ews2lFpZofXd5BkCOe2I4xV9+7mn0m/DSmn
ZxL4ep/LvryEH3JuK39OUF3jPwZhXmk+VAHZHukVay1aXyhjs4eG0X+e8mlro1qx7NJ6iphrU9Bq
KUltkSiHJIlpeuyRg2PtObaVsYZv4GgQ1N/MueDV6LbAptxvVxnzEfIBYHDsk830WpdixS+gLcI/
KVRNS7yIkIO58hJpJeZgMFlS2AUQey6UA7aPn/3bio8hUdvvtjXTArqsfxJ+JNBkHDfP3O7JtzCL
UsUXPeQz/n/P60fjQ0JyxtJYYV5ig8hdZljEfM0FO6747kybk8HOczqyFP1NLroxgYySyHqlmfpx
bIC1vg2sGd1aNvsfUhirwXKlnC9pUNvJJGiy4uj4GluK0yY/Lw5OV2AGJl4VOK213GtiXaKBjQdv
jRyeWf7MwLYtFoRua0msSOffMyOBgfkra+B920I86LoFiayAdAtAqHDVwoWuvUBLENgFR1gtykoU
FGHmEQwVldPfQaPXclppznPWi75qxOgBxCBpP/6LIXhNFTNm2pEvwGXdjxXu9d6vjqKeoWGgLUss
mQgZlmkFwklqbFb0xXaA0gucgVgHgiNJKNCYQoVchyb7pejrK3hXw1u6oSpWtKKVlb2o10UxFDbN
0Et7hklfjlZOAl0Ko9ZnLj9dk4OdCrbX1v/FuH1MLvGEIMRo97oWbxm8uRzPe8dRJ4BaXmvKWUVu
GSRdHD8EykSeo6TC4xY9t9Am4t/m1HNeEtmMmlR2p1ajLMW2OGCxqCI/laL5gHhAOz9SLAkVDdA/
YAmmpE6+dvhpo3pWAok/0vLDcDqEinvJFI+bFgSbzVVxDWVUcNYf1Zo6QeEH8XVefppwZOO97jyW
GlNTvLffoom35MatF83ai9WoHucwPAkN7B8IM5qLShNl3E6cuV6qw/e45FajLxTwMPMfum00meXX
H3dwS5uWe+136M20b4cxhHG5rgmz8rb3jSSIDB+//Ww26DRHTDkd4nJMPJOGwuQW/5MuC2V4Jlvp
i2Fhp5sq+uW/qMpub4Dd6/TX2+Qi6hwo9RL3l5LbbVeXR+PIap4IaYquyDp67tf/FJgtsf07ZGUa
BoZJNhupJTNlO9Bf2EXKWkKEvwZkGxHRLXxo3UaRWMbEkr261+Dd9GLK86gDH11xJ5Akx13TOhKz
oBPYC6y2nIq4p+ZTsybE0RqPfVM+6rLO0NQ1KE2O1m4eJTS9s6MXEI29IaSiqt9ce1nNza3/6Yo0
GWIGOlKxVGHgey3gG+Rizp4ROh4i9GHBok8+Bp8lfVBaaITc6YIue6ojGKmfDEEnvCLc5MtrfR/n
PFjfbZ2dVPAhxm95Ag8NRnMs1VcSr1gFWlZ908k9XVDspduUYABpb/bRJWAkvWn7TQtp3+tp1rqx
0O5XeUl1VsrbOwEAINrovvdUS2588SPs/ZYzxEy5C3bYsoHt139Zh5Pe9cyRFa8eNBrj2DqiZkdY
x0443FFv/1EWLnwW2wedzql5DovzJh3MCjmT5D3liO+9sHoKwBCB+2m5bWpvt/AIBib32sRxyGHh
1bdXECBEIHWqXsazBkDasIcMPnPfXu1HSYvWugCivjO5Er+Wduge+jux06bMMaKq9zixAh/2XAqV
kXL0So/l7k52lkTtzYQr6yHSKyyQxuQsWBy1DJuwIwoPNIC0Uxa1vA3a/eNmW6fPwSIXN6Q6tNXf
+kt1l27RiRwx2rITKnjxz7SpzD0l9VvDm6sTYbab/S69hFW+MHUPaYcynER5j1xCM697X1WWAsJI
/KIAjo5+qkPmAA0DieW/89x6IV5UgaFS5CsD1hyzbFUOJCrdbxOuf+xHmUZW65NeIKenLe1Wi7F+
nrllSdear6ABUoA7e9PxpBJUc/S+YteD+93ETgljpby7UcHlBbSaZF0rb/W9qgDmPA85/xSiYPH8
MJbtWpBYRC1E0hNsmVAIgIVy80VRIb/XTqdctA15XtcfrSoJRG2nZ20r8OTFfK9yHmww5Kb5NazQ
Aopr8/UnJa5noSrdGH0VM8n6uhHzyS4jYfYC2HHQqki+apc6xvq2zL1kNoHL1Bk9Pm31tNLo2bNT
dz4KA6++N1DRlSoBRbhtxG70m7I1Ql10B/ytp8pzXhODyHomOZWTngcrOBk+2P08zPW0GXB2UT6X
vgcYlLxZ4z/RwqYgR8eKCdCuokyAnKnWcyv/GnRIo8UhHcCdQbvPB0oEm+d7LaixRtEyyaWYmnbM
YzSwKA7XYXdrQupoKlj/DQY6NK8DImNWDLzonTUln0vVy1+Hdgk4huYqnXP5DUdxp1MMueV6YLQw
JKIeMKUrJ/ndKS5DMSN0zyzPjvnS9+L4LQYB5DpnS32lCIBhodNYO4/EjRl8jgs3pdSdzMP89Hy5
+1IR/bmX+nwX/AzXZ0/Ycsyf4bmINX7OLRPCgGpAKBlaU6jyGNxFq7kLuogxw/Q1k4YZf2IVeheD
DPxcs+A+mGPyCJBYuw6jadjlS0zfsYt2e9/7kTURttANk9nrZ1RpTcEQpKkeuMVmh/AOcI4ChMqL
PZTbaxZNGAGFvjqZMWIldpoYdpu9TeqFVrx11mV6DuCGicHTjjpBFk/awkacOPXmYLOUbbA+joGr
NYFR7dDLMbhtRtI/jNK4Y4GHPYDfMhxaiMlY8OnFJP2f5hVzWhu2c0Wah42YHmrmfsBNI4ZVaJ61
ZKC1fckOx0L0nd4N18SfUN5LtHUg/Xo2PbxyyDrfOpA/HTxBjBnYgirYEY3quhVNUPEXwyCABoOR
ZPXkgSZoJEQbJUXIgWLD9ueiCJRpDWCeaRyCJaXmhDsGugihxiAJvSBtwfciRPnLJmvzimNSoUPb
Iji5O2Aa92Xhe6hi83f7u2hX8bu4IB+A4O7MdBj8hfXqDmGAZI4joULR2vzElL0Q3MpqpqTyUKwD
jXIEodFjEUWZnNpZA7JV+AgVBa+8CukXrEm032f5R0EFrfHdfEWjPGBr9kBFDpXbOEBht+s2O4pk
jCDQ4FaIRU9jq5YLuv88WiuZlZa0Kwx6i2a0RMVM82eIHmK2NtvAT9SbdT2K3u25QDXdF4AgdCn6
D9oR9izAj+YuWqG1LFYCzBYG2CNXEzHu5UcmducZkKrwCsbv11CEsT66715Cyy1xPFU3Cf5Nhdwd
jq/InJVKmeIP/KrbNUfvTFsGY1sX/gogvRpv0g3lO+4CLtH4uEbd+PvgEXPFzrplH9nGSc8e4kwb
sbxe272bg4adMdjKymnUe5nDCCOPvnfGIQIADe3Eq3+e+A3PwKzinfi2ZrYayoVDG7sxSTxJk5PQ
1o8JF218/zcJOemb08udfSbnOTYYLK5Kic5b2aF6/uTGbIAnboV+gtHdaZWbgezNwUMVRQiS69Wf
U/fCJzJKHmtyT9fGyfOyEbKVXNl0akiR8C+49l1h3oVjYtNWXVz6oFBX9993euW+1/UX/P9Fu7Qy
M/vUXKNYdVg76jEKH51VPp3frx8NgtacBPwNNg6p3F0U329/e1bPxmzu0WB8wcb21KvtJTPiG1Uf
wcDZQMG9R3cou57yCA90Wo2vvqwPRDuciw0s3AIjTFH8UAFwzFhDt7icc23jP2D0lF7yk59phESz
KPhn59hbC4ODjFpUq9Fsxqeh9UmORteLn0FUsLiaajqaH9S6DPd80gXnbWcZKukb2G3cDDzCmzoh
H6XzQcNfz1AUrpjnOP4rgBNMsWcWnL5WH54ZzXPE68k68Jgbj6oQlK/mNzQ/U4JcF3JGnrWL9bzk
1EC7n1H1TV7yOR64il2zAadvZh65k+L0i0pA/+U5nyS0MUN+D9/ZI2eaJFCiEmNaYYKZdtyEOPrW
6S7flM9rU6+s0zBTxGr0DC0LqaZbOiyUf/3CpWVyqkkoXj/Bxe4beQepmKtgBVDtsTUhubJcqCvy
GyZVEuFdLGwRdE0P7Z2qjlCblRkshxVYuOlaaZcNwk6ghFdufeoQ/abtmoGEMcQHBrqtigRJV1mH
ISY7cVVWbJLKu01vfvnWXDv7Mb5kpuHHEEvaGvupPQ0c7xL0FKHMOF5bmS2rAj3R3YRmJyHo0nUj
DarRE2id9OKFYUrmt9isRvaNL2NRbQVzDsaJbA4AiXAhNMamIASML4xDwvUpPu1wi69IicqbVfmk
1esri3k/TTY+/6QDeL3KHP8Cj4YLD70smrHlMo7uOxAbOV1S3MTiYt5uI3dVeH6xfTUMsae9fjl9
VJOUC1TvGSS0Ul1Oa+h3eiYoyEsG51mtU0dT6BcKzmrwYG2nl4Lngn3//qC/8+aznNfXzJl5pc/S
KWlt5JXUtd0c5mSsKvMQd3V//HTRMy8dHhtYHOSLECXfw+a32eRFru6tDqQ2sHAlWbJMaJOV0Woj
QFDCiFEZbNiTixs8vYzNsboTHDZuIO/KeCg/ZshhWYIBBoh3dEF1qrCpW4XU+ATiDG9N54APEmc3
egYHS5nrbDZWRjimpLKvG/mYz4/ed9hhHoC3rdJlFR0rMY7Sd74FV6cegNVQzY4+rH7W5wpFBaNt
D8lnSsvkHwnthn88dLNCfxLTUnZpuy4T3lzsqON0iwQUcsi4ttYZ0DhAtqX1b5vEGjRkSetla5Qm
02o3P6C9chOTeHmhqpNTSkp0HH5qv2tOQbhIocsQIGVuz0egvzNbvPQeSx79CR2Um8rjYSvA9yjd
p3+Kv3hL44dnA3bxH9hQiFE01AQKh0Af4KTCXse2C0rv9wpAK7aFfub97sKZL0vAt6Up/CAhjYpC
35r6RI2Ph6R6MLfF8u4TRoqzKuF+qEJj5leOkExS+Hjdl0FgWS93M5a+jnkB/jol7ljTlwM1chX4
bq1QkYRFXur/zQ04BeL7ePJSelunUT2f/x2DZdOxu+sZJNH2R8i7cK3TtEPP/rtpQP3Y92m7sI26
d4OoatvsPwAgQovGPvYsxqzBwMd1dPoXS2aVjYInFjhXaIgrMcz+i2xr2RDmKCwLiAzJFQFCFnmH
CjU55VUxPOTZIj8F/UVzNRaQDQLz6efSXsu1rsKWbnMF4FAowcugoosW8eNOriJfd+B6N4fDNjHl
qaeLRlWD6Hfq9UCF42tsppjNT128mTp5iyhm6WITqA7PnY1jsGJLthagVj7GVuDKA1nfjrDJkgEs
EbvrHzxK3TZtoMsfymaaBLEN2ErSf2wPQxXbQnEzsG2wGEHinGkS4cyqZ++wyAKlLvukHcpCXlJw
XAEdLTWnUCuf4qTxkkyM/ahG4PYnbgyhkCL5RRvPgEJyXQfhZe1HyKeEVcK8YuGAus2Sl4ibkh6x
IzWc3k+z39wTjYp+OY8nSclEiNHMlHYPw1EZFy7b3hA0oDCQoTO2ozQcQHi00JWHAzDzG0ShA+ni
DCA0dy0agAfh7O2raFieBO45vT0vvbA6nRLTMJZolXxV+xfLlBeZrN3LJZVBCEzeM/pDtjmxgoDm
Yu9nuPkpq+/URKrsORP81NhWOXDQSPEups9w1r9chSl0tCe7E3eemnEhFbk2efjOg9Gk7nMQlzBY
i5GSgCuEJLg5ButDL/jzwSiggJfnqIaE3YSqX5csRBfy7srk26OMUjVYGPUJXic/MzA1i2WoW3Yy
ds7y/EOPpaPGSX+2B6zQL7r6hURHHJJkM+EoX2z22jOBvCA+jmIR8AQytm3hCymdojkhkBFjp277
hLspiD/FQ8FpSwnrnfZvPwWqTm0OA/SU0HIbreZ7bVMTbaS4RzvcXC5GXDPGGvCijSDEjDpXwULi
nvB0jAjULXEpgl9AP61NveuC4/KnPswfS0Hxs2c4sZFAjKVc9TFQazORYCSnBVNlZ7CZ1q/LtC8+
akkvt2dKuZ7tMTDaaY7P4N3glKVLiQD+OLZ4hA2CR3OTptF2I2UALwCavHU3E7PWpQREvtWaFer8
7k1hjIIIzN7/fLbLvqhcP51UgLomBgeht3td0Xo2e6beGhqkb/CPUsDCbpJVyNXntdsXUIjyvDyx
zwrnpVeJUTvBOUMFe3iUoepjD3Wn+QNzrbIDRPuApcs2H2kKHxgT4bV8pvExzzvESUn+5DB+byNe
wClT1mEirdOwRPvMX4kxV54CederQKAI+bX+g+ezIToVAtiEGJXMERuY6xHgNmJOkxUgMlHhTg5j
oU7yhM186kVMk4729fudGoIzCUKKwDP584EBOARDMUD1B01gB6IbctDZtbt68v1S6P86IfYFHPRi
V1XjCnyyBlxaIEnaDRhbOgymJpX+Ic6m+Zf3hL15V09lsr8h+fR9HFRSP/ybY8X6eLTGvxwHBr3o
oooPVfwPHSeWZ7xg1625ZR1znMjwwe2Iql4XPZPkprk5YowRLtgUKZFzUnvcB5jg3Q2u7f3fnnRL
j5/Wc5SBFDdu2CJRDRG1w06mUQ1yv2iSzzqzwXsEVWR6sEuqunahnzU0RMcy8sEA7IWjtlKCUHNk
oMXQ3ooFCRDaSjM5KHasfYP4liNl/VyENCavX4yXWavqsTAfaZkXm8oWZy2gKYw4kEmrPPWlgPQ4
vUOFFXMhBhZNJnK9GUV+rwQgSdfKF5oiWAT9ooQmX07g/5iywRUcozT/D1lB0qhoP42ko62kyjK7
ulAdhLNOFsNh4s3XKOtBvTnf9FtDomngdx7+tcwRj4jwjl1O0D6yb4f0hePGxTeQk22VVGUrddWs
mNye+84uaHKFc3EYWWlqXpCHZwUCLGO000q8xox2BsoOwl7BYknIk4b3OHwyqIbE96cCZhFWkbyp
59FQcnftWRQeULztKf+pZjncvvTWblC3RaTB/PGZ7DdjsWJW2rk6AdGUcOBRKK1LNSUU5d8gR+k5
NanvYpe1CFyUkGXPlr+fQcXsO+jKG5Fd8yXa3ZOR9L3nYdou/dEYgjFwSpSJ90BrGDQRtaPQ4Zj1
E7UTw0zq1J9IF7Qz3EG1yiX27efh11eJ0nFWuOPeqJdh27LgAC/zD5Y06YM9y8v4CiiMQRb/eovR
Ic0/Tcp8ou70zPemSWL9KCRk6gHpSm5pXqOga65NySdkcC4+H9Lf9PcCvdunTGBkOMNxRyr/VgN0
S9yx9p1Si0BTj1uAHuA71GfF5rYMTWzSNkIE3imPFXmAkkcHrHRgokjbhOR/xrro2y4huITlBg0F
4NeuP1aj2NANX/jnEqQZFzgsvzV7LaccxxEPQvQNl/+S3zI79vH+OXyQURnPxldxzozzjMQHtL6O
/nOaFU5M4087c+iFUG1XQpROr+KIx5nL2JzxPETeKkZ6nBnkdXxkxS0bHMgBFfOkigFOyrtsCD6V
0Ro0X5ZMYCwsZh5LM8rGKWKbA+1397B1R5/NUrBeahZQWTkKewTyNokdB18PQCPXrMUbKL+VEGsd
NPDRT0MoprWCItRSuNoETZmJS5GIHWT84jvXE3Y9HQwsHw7XGSjwhF/Q1vUYRbN2EKBuwcYNE1nf
b9Hs3d9IaKa5c1iaJbwBIQUlIP3rCJV8x5Ajx8q0ZWODwi7pMK8zw4Qi2LTlM06UlCNn8OYf/ZpX
lyGypf2MjaltR7eRAhFoiFu/Qq3vtt1pLr+L7HE9nWJqHO6wfxNr/1AzuRNnjGLmvE6GzcQ1/HX3
5Ks3GJMS5G63tP/qWC+XRwLS/GCC7banu5pMjYGt+F83rqaUrEiLkFdAe8p5NAGqJbOd6F1521JF
K0u6Xtu7S5n6Z98qFTh5BkqB0NQOxLV2CrvFRpT4cc3qFT7fe8Xa7SFu0Sba1TXnrOdwjzw6Q2Jp
sfwzJW9qqotyl9wINlcrIhRABouZjZ4Xfux5zsArjImu0O7DU/xF1pCN7TKFpN9XlS+QZrOcD0jg
TyC5nA2zXgBLcnIU1KxNhLH2e47vBWI+p0CU8uDEgBijPe4T/Z9kvAUSF7NuF5zpgLl7l8A63BkI
FOiyUroU1x691NQ5/CCJxpnO4+/nnzS8E59VPP2NmrTi86fne2U5Rt3nEY410Kq/MlTXEqIwhMaZ
QTYbsqlJm1fR92Fky3OZnI1rvmBtB5ZVsp41fB4CPbKB+TCT5bav4tis3lfFEvy+9tRb6O+VuVhx
9eOsZACOSI/XACB1yaz6CZ+AYlQWuRkcMnJV+LSuJoSdpU5YLGd1jSOub8ixe4hzSfU4jEUwOmjJ
af+FdIi889JgrHZcJflCxTnxOYbOrr6Dd+wo1NW0Zz4f3sEH6Ruaqj6FnDvN5DC3SQ/PZ0HD8FRf
99AdJfI3a3UJpMhzi3XiI0yZ5xgxOb5xAn1lO9AKBWZOUg+SGoJbjyWXKShTCMpvv4y6aVsGi9f4
n4JXZ62YrGT9HvjoOjUXEmXFPWKPGKKb9HvHjCsE5DRMlA78uCJP58Sm8Q4n1+A5Bl8CJx/uTj2p
A96RWZ1xvPvTf6JMpeCKDJeE9r3533+xzraCPqGptyCNRBp5bug/ptnoxAhe1dsPaKPxegjiqwgG
05eh3rUYGDEJwIkL0uxESLm6UrLgj4PYVpcJ0dKRyVGhsCasDoCFCujUVAAN96gZL/9G42xQkQeQ
laxptilZl+vqW4IEAvI1lP76+mhWrrGc2Iqzh+JVBrx/is1D/G2mkncfv6RLBfmupTTtOLQTkFkm
O+OGx3APExn97ftF2seVv4ueniBjcgDDFa8XCT6Mika7rUqv0iNgFAtbg5AfAQKEY/UDb7z5D+EE
5fZktU1oJqKOfUOblOjS5Rr2tXwJ7iYg5JB4x90oMidBwlDRDCj5qviyMRCqPmjgPuYSeaM9HjKf
brmiA22ZwObQ5pANyi2wQw8asGQ1mTITn0+cUaHOjdvZQOJhjlDvVTe+0sxFvba3IUitN92VCsxN
cTLl+BeaU5AOVxVrJiUM5sRlHfaa7RCDsDaYjdEvlQ2L5NxwIy9Me7T4QJRfnq+RsGV4c1zs28td
BnEzJRmJGusJY5FbQ3mGMy2S8ZWa9444mnKZHifG15M3fK9ojrT1MEkt5TOmRmL27xLMIdEz9/3O
rAFNzqcfhDQpdDkNXV0zEai1igmcF5ptsMStNeqY8pSE3j7ITZ+LVRvnHFPnu1EKwkeFWJUp4E5i
lN+PsoJZTFGLjzMCAtd2ABZHS9D9zI6k0N7/WV8wowH9WEY7e1AMiqBtvWfJMPQOwXzWgHcDYA3O
N+VDHlZ0BS27SGdpjoY6eRrsHi2SveHc+C/O8Rh6hcO/8w2Xu5/28FEJ8eeu20Ck8WVr+u9iR5NX
YFH6h7pz86NQnotvE0eK3VMBOTVrVBwhsLgECk8sbAFTZ/An6zfRR4CDbOH9FFfLB708nq6TZFZp
7gA9e6k/bTboibjPCtTDRLqyud/q2KeV/VGja9r5+379ZZAv0PYdSIeAH6pGQU0IF+eujSSaefU7
qwdsuihNyIEJeCicRUs7AOkLMHvR43Fm2S7etJzVztRbAb2v2MqSU6qMuLrJtvbxVXku0nwtlXHi
b5gJdsrtJ6iY0tfDdFgRFXYaXgMK+SQjmJ9uPwofgroZOkK/7nUK1yAbJa5tgUQvYrd1cZrQGoNL
RQjODyMkBYdNTULK7Ec2oKJ2HebCUbqSMNsfCQ4z1Etbl5WQRcfDITanoD6YuuzjUNX4OOmP6UQq
Jd1JHCQhnaL7B+A7TblStYvihQHROUoqdgepHRmi/P+syNxL2F5DZJkXF70WvctplZ8p6o7O36Yc
E3sF+0lMWR/aJiMArPs3qdF5e3MQ02wwqO6OD3yGeHzzvHfYf4LbbrGSghbDyacDftuPyVROp3GQ
VN2gvvqNUIpqh39VDBUnryz/cXblZIlIstmGB/my84e680UvZmlB7q9XeR6AC4umRP7ZfFZCeyJv
IsY3hK7H4b02MxeRp42RhHvbnzPHYFCI10u7Fm8SROR5BnPHV6gtLkw/QbfRiY9YBuU8NFxSW2IT
yT6q1RLrhKztUKerE8DnjKJ25qn97Fojcre/EOsNEVkH/+XV86q1eKQ57ptWWazlQg7v5qO9tPhD
ZIORnFVKQYFMLsVd1Gviu2i4ku5/UFYrWU/WWXwLD8icUweAiuk+L7RDfVUorwkthnj1+oaWFMgz
31HeYXaineWJ8VtXG3+4SVOpn7Aseqc5dqEOGshe+T4MCWkQn+x/7gCmuueqTVIQ7DGeo0AKhgZI
66fgEPAfZntKkp4D8uBbqcmdeKAUK/Siwxq4a68cU2wUHu2x8y8z043VG0sFzuPSbUNz+/mKHV36
LaEuZxZAlSx1zYoB6BF0i7EZLfQCbhOtUswSWxz1e/cMuJsaHFaK31sokoJvQTj9WB7QbFqdue8q
cdHXQyQj8GSxjJB9lWYbQaDpv4tMzGGbUKPjj3aah4Lm3YFeqjfAKq6gGK0nDWqOetxs5GM+nawS
HIOLSo6kRoiDuGVF2wPCmpIObJM13d3GzgPfbzXxNk6JZ89ZLPJQC08dunE+c0/9aV8bR/zMWkJX
mEHxP+plM2rPcrdArNeZ5prygz0Pbz/8+QiipGHryYXfkMmV+0iTWRKMQltMhs3xLf4CQnB1buZd
9ID8+rC9QbRwiGIjp7iyLxyeq3FMSBuq/zNNaBHrb+m0Yv0TPkLei6QQcRIcEVlbqaKEDbrI1Vge
R98XAkUQc3Fixrwe5eVYo0OiTGnkq8JMP0db6mcGLJEoqI4CyDX4gR80c0POaO8toSGlLJQhfJf9
aOHh3+2HA8a1k10ZCEtG7mOkHtbWhYeAr1UuysBGXZS2spBtVRzPrq8w4cVx+Np540RxDefsKDew
eQNTK1j58FZI0wxKwhooVSfX5XKsljcRbbeo2Hryu42sueWIfByYOP4AFDBCnI78HgxjaLJiST9I
EUIAS2D29ywES+k9QzTiW6tnYD/CelXue5CoweMoJnnXkCZ7+0LyV20hEl4tEQWWXLUesqzOsNB2
babeuMnvgK3lp55LVGzYH+atGvwoYJAS9IdEky1XnuFoT4JlhTPrNYMwisMxqc2Di7ekOTWH/mHn
H2MQnOX5LO0Pp4eQr/AVJZgF2KfZCnUt7bnyw7aXSlE5QPFUVXHcTQ6bT7Slo3aGSElW2T1n3xxV
E4OLkQsnPoKpyP5AJ8LOzbTV8tatzi3EFo7OK2qmZc1piCB/ssC3lNYAXe+UemIW0VlArQGBMn1D
qegaYWav56MHmuigIdWlm8RK1PeaXM17pfhpPbmXsdWWldimFBN/GdNv+k9/zC6/yNhtb2IW9+7X
BpbvEowfVHebAXA/YBnOJEozmuqu2741CN3XyB7Bi8bxxlGW7g4zPnlGmtPOcfRPVvFRApa52Ouq
t3qDZSK9C1eAcIxSghlC+GSmDSZTaZQ9modeKk0S6xMt6U5mIk6TX3ZAKzWGhv8F80higXSLDElN
ogOt4tMvN4m22CL5A6BnfwuY4H4oAtqL49Kd6mJ6wXyL5a9kDY+QX6Wxb8sTewZ6XJjEu+P9DlWJ
Ni2queH81h3wlXxe/CbddzA8PalcVwmyXp8F4VycwTRLFuHtpXRcdJiy8t3MOuYdA+IKXkGpBiq2
AC3n1gSfbecb4EKFp7es20iy6MtYrNE4guwsCIW25HekgQ4H4wQn2oXJNC6RmSg0OYSKUUQyihcL
DgMhMvViMgNLl9O5eHGT0T4m+fH75XOQpFPtxHCQidSE5G90la7ALH1iQ/1dNpD5XpHhDfSKHGpR
WaM1pJgviiLawPe0FQaSKYyOM9pa9VQhlZBGkxZegfjQEQCZOszDcHNEiNrz0n2c/vqDJ9mdY3Ph
PNwnJUFZK7u3OcW7Oo/DsyTnxDvSDoyQCTcMGnoHmYp2jl4vLj5Tl7NoSoHy+B1wb0zWW1I5RSPz
1SFWsB/rLYW29gOezPg8WJ+YcGpLDDJ7XVEDKo35ZqnYuA6S0tmRM+4J4W1Rz/rS4CvfC78yTVKq
swBvdbIgsOWEghd6vWuxGXGve5F4B7Ri28BcyyPS4ogLR3OJy/DEyRhMMQb6i8c3gqwJDzPsvG1+
ctrlX0w6/oivyV7Mvb33Fp7zqZACcZWTD8ffl/AAWCzCutU1cOBmZssybqsTKXyPE2oYUdVHmiLz
SgFoYcijuTe112h6aZHSdLUOmPy2Y9vPM7ul6oIxatHERDAh75qvNzazjS7UhQ4qRNiB22WZ1hh4
vaLYR+QHPivlNntSYBDjh6QkkIdlsXqluc3x2yqnwtbqW49rAT3xsSUiJ4OaeQeU8uvayIkbQwri
D66egycODOPaiZG5DG8P9VorwXX4XrvXP4SPjNYPu8fXOcPQLdKrZJM+K6f8jyR+OohPF9LpuKY1
fPb9afuf7Bs+jAmjxvuDaPO2mYWtHXrxgGNikJmg6z4aqui8TZDUrUtW/jcnK6+avp8XqJKSoZUd
zZhJIlvV3GVwwk4gb2Dax9F8d/JhXa/ZXT4aP32bk6WJkaVAW0ON445nbF6H6QYwib5lvXz7yC4p
KSwOTH3IxaTpQg0+dSgf7DxxJhdriiO1l0KmlTtyrfV24uF3Qr74pzWZfBDJUJu6lpgojJQ8phac
BZYb88HhWAE9Wnid8V4a5njhyWkC14lPiHdO2jqRMBcVCdQiehKBkneibdvvH/Sqjhyat9tLiodL
+8YrJtCNkuuVHKbRa3iQrMOpifuoiVJaKTEkyzzn0tbQMzcpZdEbYtHnKYoISN4rgNMYrb3WpZHZ
jaHC7pV0htsTfIXwJ1z/WtHeciqPjLVvAIbS1iJGh0I9QOfd6AIGMJzU25x0RILGwLfmif7TAMYi
s3LPVEryZQ/WrguFpzL88ZIXGpdqRyPl2OHG+COq5aSE63JaBWX1shX4qH9fNylLZsPFubObvnPr
OrTb+VsnYVDmfu8j+VGmg5OyJVzvER2ElWzqplw46QyTZoDTjLqPWGZsCjzV0V0yME0LI8aZqbgN
N1G/itn0FpBP8DauAtRxmAtOpx/oqpBKdEr+VZaE6K+OKZl8JfSQ+idJwjZ9qzHu1hQzWocWSHSC
FxX6zv77pktk6SYvnpKMfox2cO2MU6x2pb5izyZy9UQ68B0RkKjZkhNtQ6092FfPSN+xhlKfKGa+
XqFk9kxzgp6yWMHZABvSvB8km6YsvVCXEKCg/P+/npdq6Cp4LI3hiWCyr9fV2yyEZHLXSbu+nft1
uANwNFsZ5fsKjT1SOKuCFCbSpnoUI0+yUCKK67d81U+VzWpYH2Vg0eoa8POHTIu3Q477BHKEnY63
ZmVItNtYuZyl8RF2jggiP6z4dn2YEcj3+BcKgy7FJmrFE/uT+NQ9DsOLEE1QbrghzfnkYEvcgTkZ
ShHzChBcDvCgpvZb/3RG26Pg/rg9+gK7qSND/inKz3RlCNar4rbwYpoMmtk5l2CEPGvzPmAn6MKq
/ajdekuvevtCY7QiuI4Y0SV6nndDIeSBbmM9yARn+oHXWmTPn4/iPnne4CguBahEfEiMv8YsG0TQ
kYQxZScJGgFQEGCWGwTRMkEroDf00lgEnYWDNIqylKqVWX85mccYjMLo2vym0ZCVQwcYHFj5z47l
1Tz8zVkMC2EAQLAlcTXnNBg6zxUpbViLNbSrM41I1ym+I5R9w6AOQNFL4AWI3v8UjeTptujrBVRc
BL2b5+717wTi/GAPNhjxgRUy94olDwP6mHQdQFpH3DVmnYj7ff9pjLCFSjrpuI08jpPtqjRKc3Dz
pF59nYj6lpwSk01kQrDZ75inKHaUK81rBzCjTtempC6qtDOsWtP6S/zLLxSbnQ/4L/Wz4xcMeWaF
5z+rKQpKHqZAc1nf997/pN8g7cDXbPav0q4ht53/eAXeapBcMgLOj/UdTyWD6xoSBpN7os9SPzf8
TBiOviAr1mDm0dcCLT6TCngB04UmvJK0aSFbYeu5cZVQkXVVLZUU36SU5L499xu/8iLS57yJfivg
gLeWlud1yhKwDiJf0KsvxLbpctAzMTzcs5bbiTzq9XhVmG9azQGXiD4FyOPx3GOGxE08N2/MNfUN
RSRsGtvchOJaR+oJvnRqlvAM44uKnp5XqFxJMRQCr/d9bF8UTZhSXctg+zpA6Bxihx91eVqLy23b
G++pT6Px32H+qsNHtu7/Bpuup63MP5zXyyqAVd8fBGtQkkc12QtFpwROz0uHn5CMl0XLti+/uuXX
JlAnP7eX/b623mjlrtjuR9s6HMIlgimsHfvOb9jHUbyr0ioC/b29C/tSaTpUEr8IIUO8fOZP1rZx
Bp+usmySm73lJArAruI6DgzRG/tMR97kLqNpUAKflgnkKWVwqFED6NVx9yLUHsCrqabo+HTf/1A7
ZX/zW0hiyfVQnZWr/4YK4h2TFnmGCk/n/qq28JxYyVwbkLyu/plSuCzehOA7ZvDFKhG9UIR4h/QT
nCxTmHDosq8yMhk7QcNOaF/edGizX/UK4SohU8mAhWvKAYrgT5biQwSNGWDbYdDe+qVzTilkg5Ct
wAKVTFqE/oXuMM4OWSlaKw83yhduK8YNjms329qfG+KLjsbZdAV3vmKJZs6EZX//MTrnT/Brrbtx
+iN2ggyixShbIWabXBL9vXiYuO0OtklRVk21Rdtw42jNW1UFru0JHNVLP2zvmzJ6yOaKNu4DK/El
F+wGms0orFnHyzZCGWkievuSV6J8oR8k9sGrsJ3R5Gyuiv6xMHhgG8/NSkmHjb+lRrcqaZRuANpA
FOpWvkSEMsR+7yOidz5RlNRS20VmjzMPZDZ8gBZAPgLdXKW/65wLKe1MLNyUhSyo2Ni26gHiLfwG
vkESdWk3aYdD+yPK9qF4e+I68sdRuMoU6Qm7byFrp11wKEjkKUJkNz6bHDR6JqTo8gS/sOosRd1W
J8GizFA77vAh+g7bY0wcqqYjdDxlUi6ve+S68VfkwPZJJVXtvSC3PLOkQQeQQ8NsYXOD4Qg01S/Q
UqSEa7Pdk7t9BOoD/PgJoW2P/ExXxDq/K1SMumqtWi+Z2osfQyoBWlbguw1YhlbMNVcGNxo4A6Dk
4zPZhng6ERvNYUtHk/kh7r7Z/tk8leiv98o/bnOC6VAltWFNE7sHFzJEKWTVdOmAkLNPLFBw6wWk
pGlAyHPpNImT0oW1v5JbKPhPwOwEHXhdKSMxBbYbb19rja1JxOOqJA95Vt9iJnuAyFz81LOnZLaq
TxJc0p3PYWKYfEpttXR/A8FnroGD8EGbWso42ifeKwhby4shM2uXx1J9DOdwaHQ2GzzFuaWWCkrf
OpYL9pNmOqhYmBCySedns5v1wKZB7ZgeGPG9OGy245UDyjforgimGlZVasVpXGULQqNIGniFmbnC
YvCwXF3bQA6a+Vl7UGjqIMKV4QcT9wKlfjBK5TUZi29aZ4fhGX/3gjkaCWNgRW+sFubJSQBPdfgo
9dLxDCMJdaN5E9dYKCn2BxIXzzJq1NgHPGXKaUF/lslRcOPuPkWTk3I04DlqyvRjrCYwWwZR+8b0
deFtM1ARnm6CQLMxWWAd98wv2tx5fVkoL76XFT87UJE17U/+iUg1PG8UnsoE4OihKsKeczKjBwrT
jAd2Zxr5dBbUafN/xlsf78q5NurhAcucIH6NXxvyChPTxAMtSOsOJY58SWYIxSse/e8HWq+rTBth
fIJRJ9lETjoRGWuUkWP0skHghSXrDBvwyyznEi2yj4OmiSih9C5ttZWOQ3LlFLejxUVlk93DcUQl
tYZVJncOX3gxSZJaxzXGSCInUNWkAew7pOEuKTStv7E9I/nubWxhxS0A9lOYCbHp4gElJWToMNy0
XKoWnw6OUalzfWHhz9shGMPgrDL6VNXApF+WXnt9erBXPNTaC4UZJ3fNRnEUzhc7vAsD8bTJTNSF
RG3qF8Cta2uTiI/EY7Zde5N+Z2ii06coinjdqA7i+B9GkwVkVpfRCjS7Uf9EIuKvbcOyyJjhz1Nm
f4v583CV6IY5/Gm0ByoYRdJSFiRt8ZLmiwAvHVelJ+Ou9c/EbxOD6cKBgfoyagg4UPNLcmQqCrgw
qji0VGcuxtEd85xQKyPRn8ndmhEybixP2YpMQO91qwPPo03Yo3KYEF2T4xwENeUw+mawt3HD7Jc/
p0mDrw4FV0fi32xOF2+OEimAF78Xks3pH6rNDamCiZAADyKHoFwF9/DPOxEdMK+URDNbqTwNEv2V
eDygJJtVKOpsLF5nktmSGVFfpMwyZJuaiG5G2arlrG5HwgSx2usch8ouc4LCaQllTBFu8IKuYMOA
4juLx54dNf0PHiBUjBky1tMVSiEMuxZGE7yLLs00+R5275jqs6wkgidVuZs0ix+u6zshfb2mt7d1
YKwVvs1Tm0zg/lhhtDoSKbEUYgl7WVc+ET30ry8ZFRffU0SN/b2DRQ0uQcAU1WqnjhHz5Lvmc4IX
xYsFxjuPdRL9LysyPxgOoEtqB/qfL8Fuycnd/CMFXMo4SH1ArKH/DrrXiz/tU7+IkNtYYEcCp5aB
yjsFAW9FM0/mEaEduQBtLB5n4EyZmAU7z01j/Vgjz7YkPFnG7haGChqdF851cHoVjpJ6Pv8CyAPM
69xX0AGf26XGDUhPYOg0sOpczgwVM3Wmdw/G7abb9IgV/Odwntm7Kz9U2wkkQ2yhRnF9siOp2VQS
r/oOoUNvsqWrAwRwmzDEvrXcNugBRNLZYg1Xu7O1Uw/8gSW/MLboUE+SxAaA8XEEsh8SK6X7iyGK
JRrmXP4zqT4/21kL06U9ctKhDndDqnXdkTgWtXhUUxWCqewIt7broLqi+X/Y5yu2WQb2gQVmNdYs
T69RXcgIgUh3YxobN4iqdFbNqRD08AFfj7cgDiXATpEO3Av8MolYpRePc0IPGIsG8o4Cpy4DPk39
eYbejOuhheixb10qLcoG0xzyZiDlJUEA/FBx16ehNkjrGB6H8i5wNli6BPRJ0q192t7N+i65Ilo0
vQTBSAA6bfOaPRuJW3kTZ5Et8Yqcksq4tppaKPlvupjOyeUKaKRV0lkuhpFesT92xnlLw4C1otk2
z6sKjwTFP+9hsN0UzQ0EBCuZJou2wpD6rrNiqiDexCJ+T8JCaXXuG4JfepkUlulsMn41mAEO8pmF
Us78SACFG3xkBGo9Z2ooPbAPJpgYKjnDe2n4jgee1+ODw8jogP4Cf+Ym+fZBTV/6qEi7VXxsVrqP
P5lwKqPPEo/ry/pFx4KbXXNMbA1rBualBBhhzVHLEkOFaeSvYjwtzQLt9wOupc+BCU9Mu6Wy9Ht5
Hv8Pn2ABcFylS9v+9HJ5IIQumbDz0cz747VvpqC+iwYFAl/FPiVPBRs3ydOU+SPWh4P2rwvyJnf2
mdPhGelpJ/Phin0FcK6x9edA7OTncsU6M0ClUYu7kByiIgZQdM2r2f+vQG45meMCgmmZ+Og7Q9Yy
dUdrQ2vevgP2PK3zx3zXtFJVXksSC4cwCCE1L9QKebNFp/H1pwLORrc7MZ8EYn0NTF1gzDdU5Ils
KnW/iMUMi7ZqoR9AGOJZ3REsLwvmmfiWl3FVLlgb9rs3ScNu4OU6oM19YoBb3Yn4mzBAPF1DdCrd
Ah4leAjgrzquw54RMuUA9mEelow/8I8INpskM0SPpG4T1sls/7MR6Yjt+KmYGqkpt7U/CGxY977n
GWrHn5D0RlsaBQfRNyPoiOxozAH6TY8qtfV9oZtGfXgOXaoOq39frmjmGag67tcfuj4pCYhz6xA+
emaSQWennQxiy0211f6udbjaOUgNf23tZQvk+XtKUDoF4+XC3XSGNY2UaE36UxjHYc5ZdJzDRajM
tOMrGlSSUYS7km+i8/++H5SrU0JrleTe/AoIYX0uKGc1M8l01JC3VoKZBBCAUE76PKBMIUCW+xF3
NUhrxJTaWkmEr5TxmMKRpKKRiN1yqErXzwFEqi+oHqC/lQ5SZ1/LcvvxytwH9PRZs+IQGkPT+oo6
WCz7tDN7Dm6hEb5PrB92u+coKgwgLLF1IQSBLq68N7nHr9FxEcMAyLWRWOhHzgyOXltqHUdgq2jg
uGAV4DfKxphXHTjSWx7neXntMS33Ms1XlcGAaysNguyeMsyEKg90JS7M5bww0PfZMWoFjzpEJhvu
i38LtcGR7B/mepoirJfuTXqnCewlESzfLyuWjh9zSuHjh+fi8wDVaMrBgbnWS2tUNkkHmzWyMYlT
1b3j3bF1u5K6qhjJAYalb70mmRAHwBtWkRQkciRO3+gPGGNVVw88nO9zTU9k7euA8SidhqY0CV9U
/L5zv8OIMCd7izzBbVB0H0x6MKhg54AVKJjXYiIRiOA0YZRB0pX0E5uFwBTVAiBBbE0CybaI68jf
l91v566k33O54la6I01csYYRD8oIz1lQXNTOdH9Ugu+VqYZELHXjrpECRCNUnGRT+Mphi0GlJeV4
hZWpIcwdWO61aLZc3g70Fb47xrl374viidhEcXbL2BKPmv5Ff9s1xtHodcQto48ZL55p8B7QeLoG
g2SbJtGjXtoBoCAbvDCAAFojI7HOY7ZclI1qazgur/OGBbtDilLYUGnwmI88eZ9t+sp/OxtVEWPf
zeP4vE3r6/iDt90bVBmV/z92VAOq267JaDH3sDv3G3UdDzBah8ELHvY/a1458U9q6ocIFAmZTCcC
A2gFRPbWw/7XwL7Bx2xEeC41Ys6L/HSx4cOuQndmXZbVbOIy+tXxsdpUoLb7YCK2gkEJBLImgxp2
63ZJ60CDfGw+8EbyiHfMmLTD+VaEYDrzHTkD2+UWIb1IiA/IHUL4SioGOP1DAf86Y/1bSYUsO1Qa
Jcyym24UuGnouNlYH9Hv9BnA6ncv29mT7MTNLx1z1jwaQmgmixdvMZYUmhboGRdTuOc0F05mJ4od
+AyofXoaZKXtCMS41h9geP/HMbU5+ZrTVo/dOkCrcuSKbQJEg1NxkWOlRBanZ7Dqkl86raGLBuhc
YUV3jNfmnmjJEIrq0Z3U/vc/E0QhNIbSMbqoIVYiM5jRbJB6J5CpeidcqOhLPXNF3mCjOMTj1TBy
3F6JJRqgXFGLk8tYrHyrl1iqXmhgOk/Dj0rLACF8l2YeNrIwqs46YsgEJcJZu5W/MpDPLu5h0vMu
R8rP1t9yVjne/8vCZiI19qHLtfragVOIZM8n5GUwEt+9EIkU2e4ZpN1zkBMthYYXFOJOTxQBqzGk
GDTjaQXbEK/cCJ6+0Q71cYVQigZYDHUjFi41WgT5DNn1XgqN0ZsRGvUXRi8Oa2eEYrd/HA8EDuwD
4yTZ901nBWtwzhFIoMlFFkmxKB0lL6gCgKBSuxTB9aJkxnre1ldfcK2Aw5jJ6yyVk7J+y6Bmxsd4
YUjBiSaNjZBtfd+8VX0irXxMF39JlqOE8TS0/HBDMSfzgR1lwI2xDEDeKF///S2dNidKszAxW2Ds
9vB7IVtPC67nhoASKmQacJUTTvt4cQ2I8gu5EUv6Yt9yPtby+O5K7gw+O/yu5K0zMjZpY4cODYjU
n3NZPutWBaL8R7ioz0VjvYbB4F2IP7r8eA7kuMFTzDTjLDRAXegz04P0PLW086WGiUisMNz8kPd9
mneNeTRW9iMwBns+giXh1UXDDXBPA547TvHkn9lUVi8DWDq4x//r8zqR9h0ceDfyJJWYo2WaDQoE
Bc6kbgYjKJEHocyXS96HLh4KD8BmAWu/gHhTeX7xdup/dqE8tvCrOL8FHq1kX85xrOQYRC/L+hHQ
AW0ZvyLHrpk8aWK8lwG3ASdueFavEBzpf8+4w51GJTniTAfqF+a1T9v22dYNbishyAP9WutUa2Pd
nQsYbJVDBVaHI1H7KaIR+O3eQBUjnK+WLUD/riWuSFD99hl+fhq0xSX7kaw1V+PUEst82Nv34Ylw
BKdiBI+DbpaihLB2ux9P2Fqzc8gLBIUtWsR77xRmSW2GsJ/eIbS1oCTDlcGK5Oj894pZ1X7dHpEj
5N0qf+OG6iQAIIJhchhKRIk4lGknUFlJCsFHmXMonTYXflTe3KG4uEM/C6TPDk+arz33J0mlGpuC
wdSun0/r8FmFDjXEEG/b3lhEMbp+J4Q3K6RFrGlhfg4zYSE0eiE6HPnYO9piSUl4XkZOcgqgt7Bs
sD2hTU8aEY5z0xnWczO2Jlssw/lwLSfTgmIj7eN1KdyRLp1a/tzIXc3IUCzulfuBsq30+l6WmXc8
XbCwT1UrsOpXMAeA+GoU7iXSYXtU4FIcSEBsRaJJKOcoE77Al4LUMySk0b/U2lnJMkf0e5PSV/k1
8/o51HQxAp4QmM2EeANU4dFGrJOjZBT/N9Ikm0jrPCRVVDxm8mzfBorVrHHTwOYZ/YGLwWtLC81D
RjR0QP4hxQ4tSW6apRqBAZ5rjwFh7nad0qAlzc6g9ieJ+jZpdFOUEe46Q8cWPHgs1y3+f6J9hNSZ
WviaaMRKU5emd3404qJhNRNzjKD7W1vDohG1KjOJPQM6n3DgYF8lbRanGoUX8SwxSg64x6qltDKR
U77CPgcWuMyIORLRV1uOITdzY8SkqCgHgi3sAjicwBLG2SLz+pxMQ7ewerG51YAPJreyU4vOReaI
7L0/MvtaA5bDHGurFaLDzme/puOWi103wfZkwqWf5qXHRBsHU1Nc47MmHybyt/BpXCEcWvibm/rJ
bfpxClATnCLcQkdTTiWHw27KlKtuaxBWwkxtSsDd4w/2qBYlwB8VRRrigLkvHBcBUAK00leLxC5l
mWw0VFih2dH4mkOYsWobjKvGEOMDk2kXs+SSIcrwd5mkT5Ldz1BY+t5R4iu0fLpkga19z15Lqkuo
JHTghdjZ0AlX+b1cyxaakbE4E+6Qdj0qU1waUu0EZMXbH8TEnzvrlS6rVSjtLMqXN2SDnJ6Kl/0U
XpafJplebZWTtqa+B/VWpU9zrT0KuFTj+SSzTzb6KlUDMcnJ5nOswKjDAEENAMWMtukikh2FvZXD
6KJFcy5lmg6JhwxtW1qf7TBzgg2kzVuM9odXVof4UYyrUvsnnEjITR8tCPVm6LELYYt+rTrEBEmx
kO+i1HhkHJlCHU9umOjYf95K+v0H6wqKhbcjHHJYC1hJGoGzNthdmfKYD/shpKZyR9S0u797SJsr
QVpEsN33XcH6Fs6WAsJuhlUSB8HdzLZacz9MHgYrQEC3OOLvsN6nw5Dpds+3/I38ZEuWrMwEaZ02
jvNRHXLx1y+7voSIoVT5tztNMsBNrF9pMQf9M9VOCauSIZEgwn7/PC/7cmD8UM7yAbyG8IhiivuI
OANGwb6C6e6B9Xl1ZPPqY/U6A2rNbZdmHoCzRl4pVeFcQAQG637f7rm/BznDW7QPW0W+EOoRu3bY
POFp4HKS5eiNSjsxNWv9B8/asXSaNc692Fl/hUzuUGlC2y/U316FbZP6ZSd2STbiMrT+9BYqw6Tj
Ne/+iodhrn2Rtr+nc9fJ/GTOGig0zGHATiqMcHZEiYXHs/ombCyjd8yHrYEqOLxJIaSQlMXI0Lkz
3xS+t9nziGyUHKO509aiGIuEiVfUntME5pdOzXP/mw/hEc5Lj8GEvcjqFB0NX+tb+peU5CaP1gwx
NRSJ6P3HmIj+pcP73p6sHbLTMpJCfhjfz33o8Tw4a9+SEAH7JPJDN2EBtQ4WNYDjW53yRWCvOq0/
Gx6d5biAmiSZ0CohhaqVyZabWFJYpf1cVHP/4mmvL6DR6p4RujmPsgN0O36s6wqbzUJV43J9eJWw
MNSMAcZndU3ZmKbIM80d5JqlPWEnJJt3ErysEeZU8/kjfJULwxzM7QpqzbEtS2V3tq1INqhl8xe2
CrB/jJbAUkdwCNpbKsITa6HvvbDJEN8jhQKO/9m+jnRq1lBBFsU2fNQd0QEYZQdto2XVovFY1Vrm
a5EWbmsly+8HHGCPxRxgMSjifZ0hTAnbHtiiZjcphvx1pGy49S2qqzSbBUmv4uGb1PUd1OOdd5r8
+lk3fWnHtyeQ152k7Gm7o5OqU9VCnFuhEb+Y8ygTppCNR9TRi97C2ULyAagwseFF+zM6XxHbiGvY
RJz18IUnReCzisyRmFrcfOOZ2Nc2Fui9wNKusZuNDnPa3aekcmFNo6ih5wc3GdX61VrevPnsgSxt
h7K3x+9v1IpnUAP4mDNObPeD0WZ7/6UReq8eyri3aOUybqkTEA9eQ0Lcaa4yVSFEr+GjrvHNc532
6LtUyY3YnCSCpG07pD8uta0T2rRWTWXljVI/hWoHe0UQIy7LmPlpJnpiMvHLVuZyk5Q3tWm1uB/N
hs3zViQaTGObFDKd7y9OUHeYfBUjevo/9CZX1GVTrmHNsnjfE5qJGmNUzd2SgTh+dBsUHFVGwbJR
uMeSHKu6JUkIpnMICxS5Gsq/F19K1jITyfx+4a/BSKaDFNFSCoJvvh/J9NBBpBHSJyGJArpYT2HR
MRpGywQRgby1t94PhDafR3Sd95IPihrhZJXE6HpNHp8k/YNUFypqChbhnZQw04Kta90tDcKWiobs
GxAu0fV19M9j6QKCY/VO7U5oXuvJyMwYmJCKNyKuMEvOs9T/8V4CPEO58CgZQaE1iUE8Ti7I2uHi
mG0fXiFaMMrl5YfkHOoyqpCh0NFK46eNyKGQY+F8l4lRxhOxLeixHbF6GxZEVK/YPj2wmZceX6M+
WfeAafO97Fho4sTyNAhh0rLlB8GgL/ZjDG79B/+LNis1zf5OTN4Go4henRTzQBTfsUB/7Wk5iK3J
nme62aAAmFEimRUpL+xuUirITtuqWwSYmD2oarsqU3K6vnqgBUMKEIu3Y59RBcbQkCBPlJtbXJ39
UW3NoUHkBF99iMIjanBuNCzEkZ21VA0rJwC0SmYMifXL4wzKlQSkB4Yk+2+Bk1wnHZMvgx0LPIDp
v1ZDeRqvtb9DZWFkhTKM26RR1640JEaRPPnmuqRsUuqjdPa8pS2E4rcy62aZ7AaXPv5U2gyJX4Jo
sCXMQbwVjwupfveQyJwhdsLQ9UBApmeX1Exu3fLmLiEq1eJ45OqUkOvF/j9+3bx4WB39iAoByD0P
xEfrB3J4F3sQg3f91QfN4Z2Dg/uo+M9NKVG7MEhYBvXB/MVn6UpZgZaZm6hrhP65f9JPwuxmqSkZ
lqh7vii1rZNcu0Pc/L0BTTl0jGbzUfDOSazYIArJyExkB1u46Wo2i7qKYFXMnOy5qButUxsFrVvk
AZgKSoThudEg8mQf2Cb9rQGOLqMU8d+l62JetCiw/RebZiR1emsKFweTUXyWOeGGbR2djPFuJRIQ
STO9Or4baaBsD2BI9Elf1e27oo6iWBe58fJHvZ/KxyQCoYifRKnNfFy4DjCpBg0cVNkH6+NRMyvk
/0Y8Bh9m5NSVD+xJfG7MxooTogAxA40H7nP/m8ORSdj4NGvUF7AEjXJKsvo8QwOSeqSDZYnVF3gP
dSjHOffQ6rZ7WKOTsO4xVocS6KVGNDGAGiQYbx9FzmaBVVdzalZTh7QgXHFxu37i5DPBoXr36SI9
dZ+AAvoYwZEoAt5O5d2fA8qlVP0MiuNQRCSJVotiEzhkLCaE4fPxMDAmbMgGYcAYUJNzfgCkzgjg
xVLHrGC7heKltgOEta99MrYxX2I0h0arUbKADUGAc8DJZK5fuL1qx2u3WJMI+rPhvNYrZjGI3yZf
WO/ehESbtHsQiBa4NbWo1wC4S0RjsT11XgpFcGy8mRLwb17o9bCv2hMQZ8D6RNi6aPXLSo8sPaBj
gxAJ7mEYLQD9nL6EBpwouQu9QfRx8g1CL0TZe3HL6TSL/4QSlFKaDO33dp8oJtpJJrOMdqSd6uwQ
j5AKhC3vsZxKJQY0nKOydY0o42oU1j0XOlDn4fg2ix2H6m8HGtOdgbpPJevEcgfCzBLe4g6XQJYv
oY9AQRgEfYsV+hmQDiNoWWxxTGXdX1RCJlYDz72uYMBnV+lrJ6LOsfaEG/qDQCd+PuxJ3KK7ZPn7
O4ZYFaA7C6LhE223Knao26nk7Qf7+RRpU4dMY6P0hHshk9F5eBEsJstTdrYw0eqY15ure0hcXbk5
yNXTEbbqQj5PLMWm24E40q7q3BtOy4m11oHpW12WuPX+uME+NTu4kf5p+kGQsE5GX8dlcnGpyg/Q
uAVImU/L+BykAJn1Lwnc4w3i/rjfuZODqu4Lvg11M6R5VJTZypFSEPjueCyaEBZOMDJ+uKlIqsL+
2FXjV0cEn6FVw6tsgHTWFh127+HUmMGOF/5+fALdHiVnccTyZcdtwDUemA7TS3JwHurw40OwzWRt
SgjYkfejglsu1LFULWfC5ac17ae1h7nvDKulE2fvw42imsFw7E60+8lOvh601qTuBiNPKFx+0BlN
NFfUvVeUBr/6b+Dvsyr2gq5mVjO2JaT1wc4GShcD3Afk00GLdesXUcAZJ50jsUA3IQDI5wdylBOi
txqMvKIFz5zwtH6bABvSifpnpHZ7tmf8gDe+Lgc7po+JD9oKFUCtq4ZxsdPl+EtPjEpkARzS4lts
AdaUyzhkDN87rY4z14jGSCwjTmIdZC14SFSq9hxEp7ooVWBoAHa4UbcczR+SqVWSGpmR05M2fHGs
AQUVnUy5Wzn21imlOo5mkDXO2ghMxnqcgYnwpYJCeciv7vFq9jkVuUeyEbLRhlek3TEO2eNHpdKv
mFBXapqCYINKBUrjt3Jajnbf4Mww8kQq5bw5aoiIaakDpqjkllvxXzZ3Qn2DVAsnsZk0eR8LrYOH
CitGFpXnStyFGlipqJ5prJJxTFFOWfXaBVCLkLwtoNq8jMavAGf/bR5Gi4ejj3jgICP7VrboPHST
pxJLo8bUINJv50laIh3NH5DZJ2in9xnaptFTrNsqcMcYLndJyVKpauZTbobWypMZWLURPSXnCLSs
5I+STQHqzxNOwD79RB4ONth0Enhq+oPdFkI0YnGUN0dxVNld193N0fqvdJH2WPmU5QZvawzJALTU
/L4a/9r8BqzrZVRIjiwZ54ULs5rzQtnCl0sAGPW3Rnttg8cd4hIub2NBWak9JTBfFAqH1SR+ANaT
rDkIjMunVKERUDlXfNG4vOIn2w1ce7hapslfGsDJPTR1TEOVnK+ZtFaU6yhcEtXA+rfycu+C7wGK
eaYRFDolNA6uYPVO4eA/TfJ03CPtf3HWBd/Ow3ETUsiCkjlz1IQvoPMzroHvr1FY3kxCFrTisC2r
qj81ATZgkm40ebTYu9GHdTj77MijOkF7oaNm3lyaA645gD6Xhyx22rSJl6EhUiqNmofLaOpo0XCZ
1Ulbzk+E+TuehAWRvkCHO7gtmBOs8PFgaxT4Z30O5llX1BAxs+DT8e8FLKUIv4Er9nQPd/fcZqYl
5Ufn2ssZzwdVH6NHgcevpxULyNvWNPc7oVS/3RlNO4zYcv78ivn3pH+01JCzBhu+nGwhCqDJZwLJ
5/nc9SDor0pfoM3V0jFNCEa9a6evS4BuAXOBqwn7883eN1sXm1SntrvlBeDPBP3qQ4aSBDYolXDN
ATbFnQWzz2pCE4THKqmafjJhL+bok7hH7W/s9a4TFaIebEdeLsTTx5Du15s9aE2Uc4XPjL79BURF
pqRLu6ad71s5OvPh4wVAdRNr4ClpmwNl1byTwNJnH0FN4yrwQmvkhc0ED4VaOF/5PfxnAS0cQ31l
KWnTbZdn4y0sBuTeSTWJ7uWWbEy9O7GyRFNlG+Dmt3MtpMfLiEJlZpfXWzOQpD2iVW7IBqqjueE7
PBpsuzEMYI9aaMwEJJ6E+/oEWlly33CUC09BL/OA9qKv734nwBbe+ohtyyfTGUapiLbmVmFsMQZQ
1GEvPy5FL61Z++GtS2hFi6a2RcaQ/+c7bOK2nMNHmGN79XPPco9hvWBjj+q+TwWYvdWAtgUxQoq+
a38cI6sfqdlaAutlV9ct5hwvnF+wYJXh/i5g+6LI0TqNRlklOu86p1glomi4xvYtrCI7VYLYpY9h
7NtcVd1sqkusCDS45S7FZ374dkM/sDeK0jWWdR3w7a3xRSM18OhN7EPMLSBJ04EUyByrzTdJs+aw
AvpDw3/W69JLF/WFdT73sWRcnKWFNSnRsUXlZqvS+aVX5F5K7BwxcrhWpWso6cCW90PMTH5ckYmY
prkw/qsjo2DM8XjrIlyP60BeBcAEaI9SdxsOINFXNePLm1d0itfoxJ8+1Xj6H5Bj7SgIBKYALs2w
lzM9CTZ3/QfhXlcZMXiZcausaZ8Rm03d1EdFi5jfsT6FkqIiQlazzYTp51BBr+6tdeJm5StcPpYk
FeurcJC7FadOQ7C83YZHiV4LMXxuN2Nw1MyNq88No35YcZCzo+j9PTPoYd8JYqwboabgDhX03GtV
P5zqTMT/WtZAhrseD66g/pa2o/7PnZfSGfzis9H4fX5QO2Pw0m4oMHEhkT7uC8d8uTK1ey3uKRnt
QAUaGgbthe3ieGhNCb9l9dUI9nEKQXCYld6EI1/hjtPDqcqkFE3vXBsC7zyyUHK8678IvQMaT9Bd
ZdehzDVRR1472UcV6wojh7n5h5KinhG4UlwbJ5Mk7qxmI5fvUroD83sp5SmBeRk+7w25+CaV9KRo
pc+sBv5V6Ceemag5EbN8DO9wgk9J8+KV/ZO02civpFIz/15fcpXkMy0R2hJ19FmkWsMqrWC0BXx4
hyGEUH/kdVaN0NutqcXmJrrJv+5sjHXXZjHGwf9O82sPdXZ58NjOs0HlD7z2mrD8tU0vSBVdYt0L
sA3QEus20CfgFHpU/1Ih80oFCfCwbr1yQ0bpVEV63upP4leeW+9qUTEp8V2rwRC35eUNlMacmnAT
4FajF+s60snWwlKrEILsyaRoRxoH/geZ4/HZGXBuRL0UPWXatjMGEL3ZxVOXPgEBrNKa57RdT0ya
vkkhQNVWXP0U9sPQ2XGt4MDqtT5Z61arbpmf9S1twMO1Xcm7KR1p0sqz+/xfEf2Gr60GxQ2xNo4g
ArF5fL6vaCvhpSnl/mO5jKsokLZc6MtDEwE4zQngMil+gPKHfhx0kIcyOQXLV1fuAI/v6rTfoa7S
eif1FZeFtt7kDW/3hXdNP9il8Zn3ZNkM/Vy3CqZqeh4q8DbTDEDkRpACZqQUlQlOtZZKhjROEj1X
FGkKLBH5eKFMQHKfCHepuaXTOw79f3EHu4ltQIy44fOaaranOGaqaeW//IvHtcFsNOyHQOg82vHt
HQJYl+rlEsr9FgO/ux5/ojTVRKfdWMMM2e4XhlC3usoHfxWCIjdxwZUT3dafvhV7j+pkla6xnxCi
fHeG0JSjwvSMSrSBjXO5iDjBdom/jHYPBxwOwZhNSj5dSNEtGvAghdJ9+9xuzKmupp8s2nOQqmMZ
WTk4JgcuaDn/DXQNiD8viDg34HtZcZzjU7zG9p2/CgvaLPtcWfVRdWiWXvO3Xypfsh8QrDSN0t8S
802Iu7myUp7wqZ4KmCFhKsBC2oRsGfYwWBPc+hBsY+A+cg3hqok6VHjdTyPXNJiDzUfjGJoyoPCW
mclb34QYgHKxybrhTRD29F4+LfXVZ6+vK9/NnqXXv7LemACt4AmeSv3Y20FJTWQORg0b2IZIAPAs
czFm3OnK4OU3g0nm34S6HkWjGsZZmt9zdCQWaiJnFRuGHutqp0EoLir6riX9uL7l+fPjSvBWG/mK
xkh+fcIw3QqTOGI6OnuEZdGDQf42lp6BBxUp+9gJKYHk9jVGPTUemOEYgAtNxzR9KMcdWjrjcWQi
exgq80hK7XRUXGX8hCaLd4fTtktfMA8mTReiREYUePNeHKKIktOuZJvvLdMBZslagYFevUXVZcqe
Q81D2N2UJMx9s+jHO9tXJYR9DGivxA4KmrkWZdIxNT0di3128u1qTWFfWljj0w3zxgEITFnkbklB
jxOsM8igSVGhNx/oquItnjDK74dgKc4lvVWV2EO8UFNz9gH8JBdhhTk1yBNwXRQl6WYC08qS47mx
EvlTcW+GrFQgUROjfi9EM03pXejQd7DeHFrlqaLPEX813arnh6gh3OK/7PD+2bW7wopLd5TcXmbb
kKmXpOJZeEa+bnW7m9sIa/7icZDAwBmpfn290vWj0O9bgM6Qw8u+5XqKwabRMV0fuUz8w/VbP+oK
Ici/cjqF5RDJQvDn/LlD5b3fG07CZbv1E9A+o5MKDhSJksjWjFJX6YEFY4NM4ckLnygstrht4kbA
lzx0aVXX2zQZB1aS/EewCCpY5MdaWaSLREckJXKxGLXIM7CPnjUyCeMBReQLl2fPnuSm3fW6oxvk
8r2p5QImBKlxfvQuiGS7Yjg7r0Ou+VrYwVJpYNj0Mt0MPynO6F+EMI7m/DWXoGfEQK7iQQeE658z
AVe3RFbEvpw5ZyiVsrw5xd0Md+xCycuo7BbKbpaVGx7dceCQ/62nZrLvA4acmGQgU+O1NVQfwloj
DaFt2LgyzKbQMVe5zlZhO8H+wDdaE0mHxRf5l/z5QjY5uVOZ5IFLDwIyxCPovDBHEc56oErcWm6v
OViwpRFPq9Qn0UEKNy6rq9BgIw0C4xrs3PYw0QKYbP8Ym8kfbxSMuBtfMpRavNHvTMg/RFNOF2Hz
kionAX/uuPaqHbkIwco5gY30yG0eoWJNXureRiaCHjk846pfaeA4WYRGUEDi+72UQMX2yL5mKdO3
d2DhhSK3p2s85c2tDBxr3UcJ3Xhx8lD3TQdS9HsbxDvVhnhVICHGTrSHj0jPiYZGSwHhOWtoO8eS
sjrXy5o8eCW97n11bhfTDnqZVQhhFcRUybHOpdeRQEG8cK1zqS2fM9E3UucGLhe1Xj+HuC3VQIK2
B8koJvjZfVK1MbyFVH572ykvy6SsZRqxW/NSSHq/DSCd68U8LK0yj5qevTtyswWUw0+P4+W12Jsn
jruykInMi8Fm4J3cSy/Z54aqhqu+NbAQldVHMeUehF2TwhFg0P/Jv/rKeTgzMvyKe95TiVthglbP
SiZXeJSdcpkUUfTNhgSMRMl5Zwk1BqioRuS0som2z5sgy4JpcB5a1Ka3FknR9793uz2flTsmBlWr
fSQrE1KlqjSCLmJL0Z06UC0CriwthbBqL6urMx0CDn/gxysWm4AxSdGH4G5MBVCPy0QpGPI0Kbd9
SM8yc0hbwi/S2oWuudA/miDZbmbxuhb3ryZK9uQBZF62X9hBrv2gV7JdwdT2Y0Y9HSRx67Syd94d
jHcgt6Y9Lo4TJKql1noMeARUd5fq2YRY5/k5oYB9KiMOkqbhOIFEy74X3L2gRiWQHJalEpwcwFi7
CHu5VliK4j9g2ON+/c+ZswrS4dGniFM6d5JZs9mJNz30qMeC/jAodpX+Ykp3e8HZ/FxCRrIncb+y
9FGyNnwLbXdd/wG0o5726y2/SdQjpiXw9AIDFNzUPG998KzZiELbIz0e2bg62jhoFGT96lcZX1Dt
661XQ9NZrudEGIeKnW280HeX7bL1By+tLyGMCSeFQGkWPOfe7ucuDlUsxCkRzOmjMQOo7A2BIQS8
jSc91NoS03bHa486pAfVGuSncXH+hNiM+K1JKbQc03pJzOala8cCnFz23IDbGXfFkf9EetGYtfuI
Oall9NQhvd6Rn2raSWGk0kz+AIz70QaPvFUz6OD6DAAhZwMqmWBQk4xt+0wmYD2SUGTIocZGgsXx
BuT0WHdeWQalzbE4soNa5pyMycX3CQQS35ekl2qVYKRy3NiHtdeOqd+7u9KSCaoMfj4Uww2ooujc
1DO+OLw5LiLgTSODPwUAhlTr1TUASFBMFJ05t/OGImLoMtCBK8vfQTrFgdjNFzcULOgFchLPiT6a
GkakVhsVS2oABiU9rwvrfS5ZZKRv5Kk0XfE8Xbnq07tWCjDS76mK17S38xtyc41+0NG6AO99U29v
Rd97FOBvdOXXTicmfUgig8WavqyLp9Hqg5C1G+RZnLTor9xlQ3flMMnL9TRviDfOXyCBBRv7YVMX
f2AE8wy11Xf+NPWbkSk7IsD+J5pen9UDHa3XgYyZJaAzyZHW5l0jxO/oFy6h3OWhQ/h/xt/L54pm
0Rx2pL4Aw+ajkI8v7j/OFpeNCs60/o9AR1ZqblDfaooiWRo9ESDtoxOenmgK+mN7jpEmca2nky/D
3PYraAqm5KQBCzAnff/q8JnENcQS6UrzFooMRrWVIVjTktqECAO6R78kaTxzv39Keb7V7hFevFHO
xdHt8oowCTPa/cMEy+MG5BNfHVYH9r+Or0ye8Od844Ef2nGujSCre684m30QUUfZiB+ccT2J7z8b
81F23ax5JN3aKsvZc1+0phVtrlG+54Pf+zgmbXVqnl7fcnp1EYVAbbXVB1bIZs4EGy23rxobX1KG
ZOLvC42MMvMGnWnJWsKNHwkw007KpKrGr60/xs3vGWs476q104p3oUTCLAvdRvvKcee/xlJa8+aX
lbuXaRNfO+LjwWsiNRd/u515JhLcrFkX8BbFh+rqyR1D9I6j5NWfRfSpw97t+uK8rQa8zKa/Xijv
RzDLlw/LCxMqo6B60MFhbhlGFzn8VYLcpCf0wE2e3LEX/yodRq6yJ7m+lZ9OrshOTzuB4Fcp9y9F
KJdpCv9DmFiQBSGtUL3x7DF9e1e7eojEWmCjp7heBGxIgg8XSdplrbjG06+5bUFOlK7aeHyQWo+J
jBanWipmKUs5jF5ded68TX+GnUagH9MAGKwRAikzRjrfpEzmOmlUm8p+J4rkVGLMlOm1EELo03jc
08TDPXR+otqpF7699bgDK8vr+lVASI6OSbYXhydIcNd62dZeif3lT+cbw3zLmr9cY3NMi4m9GKBo
ddLYUll6Buhw4dPnXnvbFAF/hRY7GOqnNuuNEsu5HBfs8qy1Fyvwnvd3lExB2BujlRtvtNA2/TU5
n3Kh9e9y7mYcL/ZLX0LlNS9AMZv/1eCGvOIG25xVJRxQTLY0WVilK3/fl48sizx5HbwbyXp1wZ14
NgrOyheqDfiF2my4DVKPlchhCWRUifFLIlVNftViK875CD+v90QGtf2nDu2M3p1DmgLjVy75fCXx
vBSHIYeH0hR1ijS5/hsyVU98n3pLgMpw9gFeni7OUIXLGjbDHQzhiXCs4obdIsAlZnCPfAK6sDG1
95bUkF8bK7qA0Ikv6HVelIzxfAaWuM/N1vWJiCw0rLIm+F1v5LHUlf2gx3I+xBtmg9Np1/W4t3e/
FOex/GiwK91ogt0DTQHgGUd9SJCzNn4cTVEBOWFALH64g18qsY/PtPR1azdy66xnn+ykGywRK+G7
/E195ckZ9Imdzeh8RLyTGmihrzm96vIvTpURDVT4Kp0EMtbvN5d1Z8zzyqvXbUxuEXhTY4sgabE9
yHfAMfm9zx3NrGJr2o4g6ZQvVJp7f/uzuhrWtewWPljUzWQ2rmPfJLIFtCIhI/cKrK5RgXtytntU
zZS0cZdYIAY/4Qtb0JApOGKDBFMovBoHp9bza64xjtk3wmRtem9c7vxx9++EvywMyE1TZDPua+h7
NBtHz4Xf6GVZK0lXqHfglamjSrpD4xOI5LxVzZ61PmgJABQfWO5zMQWYqTE7kTPY4u4t425pFhtx
nAO+RQLOsFEYVK+YBs/0Md1ta0/tl32Mi4REfE6f7LW63HaKrSSehMCEzj7rw/ZIFSYcj769WDOz
X/iynEieZhHLINxEPzlp6O7BbKsDul7/NCbPHil0wLSFXLcE9c3NdnDys14QOLBlAvC7JHuAOC0j
Y1/RzWFZ4ZE/bb3Al6jCC60VQaTr+B81Pphrpprn13Ql+vgboj7deO8L6ruxzAdffVcdRzt1r7DU
329q6kYIz9znw/z4crHEXfZgGhYI1h7c+wQqynFt0b/awNLuUPDkrQItrT9b74UD3eac04S9UQQB
EFOdssTvxqh5Fj0zpkR2Kv0w0PWR1Kwnq2vULYKTfYPGbIQo2Ssrs8f59fHcJPwZvrTtFF5ffDvx
+GSSgLCxu2RHM7ZtirtFz0Gf8hL3jWxf7Fp0EIMGAnsaC1CzpU0KeSrHCtKI1qa+yo6Q1S2AI+Xj
FKvhxTSwLTuApiUCKoKUmKmk+NomaTuu5D0XC+sr7A5oVH4SRrdu6iZO7sFKr0tnJqJHpNybIZbt
0tWjL11MxP2MnxBhAD7ZJUEvSsjhpC05j9EOuHYVL/RVYZj0Q4+f7yXoFCBD6EOgqKDU9qzbiEvx
d1g5J5jQqA9kQtSlkkYcIT0kgfcgQZd9aE7ydnuvUfUrZN2kQuKz+YdCtTOEbttJHhOM5p0JyN4Q
jVgLs+rWrrliaSNB2fG5luPGasrATYOgPYLvTfXnZFxvBsCT8JEXmkEJBuSU5KDIGEa3bz4fI590
PZNEy5WeLy3E9JRxp3zY1173ystLqoYSeGqn4kAc4Yptf+chhDGRYRRlX5TTj4yZaXQbK8W8cuKx
LguI5KeaxeWv95CHMg1mDeXe1U9HPQu+ye7F74SCyURxkY9Cb4XFut9E1ZCJAWMXp9LpbCPZIUBl
WT1RQHZ0xwTEsgitjRziq0HkYvd/hz7Ic4QL/NfqJjRXAHuM9PCk5isqAVyEk7wrcEoFr15vi2xR
4y5blf+q6MdWSda9Ce0irDuNsoeKFyAJ46U6GhbhQ09YtXCU7eq+9qWrUvUQGX4FIqJ1koh68+tz
GexdQYzkpFBgPN72Kaz2b/Bwx8woQH5ilF44hx254VimmP+oSi2p97AHWuM57rjUJMdwOiUAPOVi
EblkwJ8GGe31eNV6XwDV3RxA38y7YKf8Y5pxD/VfE58W7Yz7kmxYBiUiayJwXGQaPw3JXJ26DKVK
ya/8cQBGbsPi3TyJ/H1hIeSFSKqtoYENkHC5IT3xDILyjeTuDxwAJEj0f5zt5ghxMjGQDgp3UciZ
U1Ksr4hIhLebqr3JvgA448I0qfogdbcTSwPzyzlDkYRuTZkP8dD7n5UCEC7OwVRad7P2wbnyMONb
7mbmXJuiVA2UF1l8YT5YYxHQ7AljdAfQiM6N6fFTE3worMyZcNkJK7A4ZnMpGdo7UVgeXFHWe4Df
6W4WUkD4gdwEIQASP0UWUdBAmajnYV9Z7a1Qs2LNBjyKAB6TrO1SqAu5EHJHxInhW3we6AUY5/CW
A8GigF02nFi+uNBEb84hO6h1qJLViZpEjfQt+uCZflWPcHuJFbpUXvSVJ3o1EhHcUIdig8l0Izey
oiOVTc9TSdr+alm6qv6mp2BlmRqeznFc6oPDa7OaGUh6lATrc+lsEq+AHzwZL+O/adRMU+v6U9BI
nuKcLPuJRMjqiglOlZujrzaTANe5biaucY5xssm/rjEOVwoUZzAwLdQqpD/SAHv/mOr3D0x22HNq
bKxaIYXxFtVfF0P/sqzOIHjk2WkPx+A5pA4UB70wyn0ZPpWq2wkGcM3MM1Ke5JjnGnEEVnjWiQvv
3srNHzVT7j0R+/jxZHnIFDDdV1dDzkbrssvnNJ+SprZexOcjGdYjI8XVIPWbalCXDqSrHhs7FVnL
A3DK3UElV447Lzmg/XqQtOhf75YXDqHhCH5a1o4dwqMx1FMtvqaxukMe7iYkr2H40QfVLm8LFiZK
BEaLb856j9eG4KbKwhyR9daX4AMWx2URfESNkRwd5ClVyU98+D39IhRBSxC1m+EBDFgYk7qMujKS
u+e3sRqDRIG2Ysym0a/Hvs+OLMZr3VQybas3pLq1x6c9zjsR95zhfa2WWrcLTOfDw5uX7UqXpB+d
6Kfcl7crDAJNKGMjTVsAAy0qTeEVnOYQ3f2ncvDtvuQMH2PihER5fF88712yXzzi3WBmXFtMU6V8
CEuEzfSRLq7GCsWxwEwr1LQYRoR4Ti4lC4fw8nB90zNi+kH3TTM/eP0YWeS166RrSnExijhstCX5
ENOjvugg8njvbxlYfcNwF1sKsCW9VR3J7brwUmQLZBDpcuFV/bIicQF3VSLDFQ2exQuZczsTYCyH
/UJuKWbl3aKl2gVPyVtH+FwneXF7NXPdw525Cv9pNuQOnaPcPafHrKfdq4Czgk0tc1xFhMvuPDnE
kQmxMRzBrYKR+G7zfX9jwuSS1x9zMe+gwCJnU0rsHPZmKk232IIAITwLDSDRP0EVtiqai/cX2MFm
ktMyywpw/G/Enr3+Exu2a7Asw9RF52gNxr3+CmiYhw4WrjpC0gzHOnSX0kRSXtHKJj84kTq3+26x
G+F6cRRWBC4P1bQZvY+YmKvEW1B7bzD+2+qyb1lC8lctCUelfbegYN60fYHQaXAsiZucS0XezfYE
MRyjb7K7lrBmsxD5GqCLMJe39ZAcNhmbRuTHrW1/LNkYGPRQz0r5J+YbLQGARkjzCXJr9BCgCUx4
8vAFInPgjIcN1q9iSHg5lKN2Cgu+IkHlUSd4XKsZwfjRi9QxyG9X/9ebcEXvWsFND4Ug0/LGtRYK
3tAjv80f7NqttNJVvw3Q38zHTkAk89CuM6AdkNcB/+fFl6wbD5JMhJImCumRjjSs1xHcneBzvF7A
VPcqAt1PexCmSoq3ZTyJR0LxpsWQmQgI9eWN3jEt6VXwSFJDPQkGlUpnwcOoECtblxCGBXbdU9T+
c7xYGbBhljCg10MnbjIDUHlne72HFLXUGMJNAMXE9n+LIMfR8zEAgZ0IwuIqRobDyv5TjDw2XkA9
Xdnv7K01lIcfMd8adn71GE4Q6eBJpLxxTYLPk1VLAOzosSwplPALoBovJ/mOnJqArP7naa78XJye
V6H9kNZgRQ+7w1tN3HVSlPg0VZnLQ8dTCx8Yy/lye4G1MozhbCYeeDJiTEUQzxUDGpQsJcrwaJVT
dbrXLqPJY3lp0odkoxXsZFgLzj1S5CZGc3fDKXg1GR4WzZYIVuWO8iW/2oxkK0BRAIQViZZ5+eHW
Q7Tw9rDsTVS7Y/CCHEMA6Wd3qgnaiXlGdLulC0QI5i7CbQ0K2Mn5sF2MhE2OI3wEIWhNKaD9Ohxe
GNkQhJigdAU6UcwF4xDe9YZKBhkGPz/DUPpOFVHI3q0hgoIdhI6u332KFGV6Qj2YRZcaIqyKrZfz
1todQcArl9CUIBKIcbrj5Nqnwq31CnNw8Yrxz3uhQYg7Xdma44plUrLGzTulz/qMlvdW+tBbs11m
29h1goUxxvwRz8WxU0Tvyv9V8+HXxLzOAOvaNz3SRt1l6WfNIjOfBQCBeX1HTLuSQ48lY1QorbsS
UBqjVeDR1XKHDRQRQql6Mx4GjyoeRNvMd4gdnl35IUliiJu8QYsaQ2N5nzjojQX6YbNrbxxKmR5r
zswgeXz2kmuV4DTP38l3jRIHD/sL1LSHRVOYPiaWyc2F0Wxu0o+41mK1e95Pv8WQ5U8Yp0YzpqdR
eqgg/B+FY976BTPP/R1DT1ScXpMzWJcDiRarpmIb8NNTpgm5+wmmGFHZtYBQbi+j/VoyqgTHdRHw
Qw8IkdTcLgWpVmUvqmm8EcgX8n7NYsBBYEoc52SwxILczTlXA82BRmxxzSzr6N30A5dKUcvhXnCy
F1/pk114AlsPiIDhyxM9WZuWcgs1IjWO6d75QkGHFCbTpHjKtHffYFwe3jLKCyaBTtVPsBVz5MvX
fZdokm9ho1gTQ/iizWPpb0FzW9usoqnCwJHD1ppT0ryhEMeOivf99bFnO0CjwKjdRboSDn7mjXQG
HF7oALYuzt2KY33vvJh8XhmmAIC7ih5i4GTuVtv54erNTJYo5LVgusWVHkutzoZ0BwletheBHGTA
jllrqZhdAFOEqUsFgFOWcGzVtvlr7gUx+lcDRj8FfYMgRk4/aPPOKVq8nWKOHKXt+acDQKVsUEZE
JYEZ0vbCv9qanbxcedmCInbiG0x8/E58lvIewjB309KILrRdNRnh0o6XCk4cceRQ96MJz5Axo9za
lhokrgIL9zkICOurOF/NibJoQTMjCuzu9OUAemG9g5hPsrG3ZZtXzusDD2bYgYu6RsV+KArUM/cb
QCkMxPTtsskU2aTdqTTMXKFTAWPETl6CnNL43YzPjjMYi0whF0lgxln5jyz6ExiOXYTmxUS2p4AP
AjrUVf+zWOU1VKuFVHivEfYjSDDPyUy6f723ewtRZEEui6IBJBvtjMa/cxlSp38JGNIJEYNdZ7p9
WM9wZuzpDkQrr1QXPCjojkitg2v1O3gtHggH4yLy9UV4Qa1hTRdFdLtghQYwQNSnK3DT+7tUmNZc
EFTr9dqbLvC5BLiQH5y6yyXeuIAClDFgYFdh/BoeTs2XKfgkFwm1E159xmsCbIIuoPJh48inzOIe
v7TSObAIDrFh4tcTTg47/ujdw1E4+w5dtFEaCVlisSw/Q6OiYSfYfSTXs00l1x8L16eZt5CTYdlr
q6KnBPibNP/HpiBzs87fKTg0y1tFCHsF0fBh8+YB7ViwjR+FLeHd4w7xWAi14UszxtyJfzrfxU2G
yvL2XWdii6rKI1GihWMmqJ83rxsSWFymH9xVbLwl1AJ2h6263dGAXIFYUeLd/Tl6DuXkolvEWBd0
z35yc8041MxvSpMGb1n1tuW1IhqQpm7JWZPBl9KBgF5agswr2RRmR9JpEbLTmmE2xesMMGQFwlH2
S6wVQGfx5kqp4OX82kV14+39ozzsDrDwL4bozBmCtki6iUGxnxLf8y1VQ/Zu8BmvFWSLJsODifEj
8syg6i0Xp/yly2mDahlDjX/TrgxCcdZBh2ETxytMIz1xwAwzMs8VRdWvQjSBqGQRyWwuj/1O/YPz
yQigyHvyBQwxYOBYtzqt6TOU0o1UxYcgHIKtNbT5rCAE+ZmtlJo/I8N5RGw5NN3QB6OsSHnbqsLD
LjcN1ZQXjrZk1vmHAroCGuFoh9vLOvLgZTwXtEf3+YFhO4Ur3CKRQF6gYyMbG2LzrMvgCCUaNwNK
rQnZwa3YLdMPUuWOJ9iISnamfUwGyyXKdC9fctPwef/WG2PwjWRHslo63pHWM0BLfdwls2V1qxfe
0fodqNwso6moOqkduOdOrzOaL4rR0jcDSrvuODojziyNcLrAXnKMOHft6W5DvyEJSTQoRXIme+Ya
z6jRVu7HbM6OdGmM1Q1N7yIQaWkCiN7oFflRo9/Zsf8O3m7+ylURkceyMYvQP8KgWKUdeWamY5HI
bXVcriqm1cXBeLDm/iBr0SfTYPSHa6JHtI8Y4s9MwCiJxoDVwPNfP7RI2YftLTfVzCf8U2sBkiVm
d4WQIUMol6nDoqCJsacHaEHppJtQyBfJ+dqcJCRLavwn8hpBkifG8rntD2JtAieHSB0PplsUCDnp
e2wBBsWcxiMQEi1SfeWairD9XFVBrFTiGKzF4ddIARF1VifM177Q7GORDCvc+sF9smHOG2yo/N3K
/FZp+j5JJsKmXVgh3oB/CRrfySIWcIgcGI/H8Iqt0iE8LlHxi5tomQsQkvgdyr/6EyOHfHIwiYvZ
eA/tsOZH3cdK0PSvV5X8Bj+N/cGj/eW7QJW2+lduzQrhXrpzBdFtjM87FhZg0nZsh0y+QidWMwbV
dH/6SQDu+MtRkNffui6A7+c1RMHU94w3epLLwIdCcCFgPBbL8hbpKsob5z2NX33r1Nqy4D+B/wY/
Ib/vmEKAjljQ1/pgp0o8EKgGTlgmGA4tdJ9+9VrIrqQ+Zn2+0UKkrQE2bUeLFrscFx0u8bycc2aC
lH2UfaooBlwWdXwXrMtvKd90shpbvFzbAKnZf+U91zHXmNK3NDebDHNSluJz4qQmwGcy2/lFPEhJ
zV/dFk0OWfPBbUYlxI36tAADpXIoTgW0IF7/M9tZ9+CFHj3wph4gSawiCEE9Y8HURP4lcYj2IEGY
2TGNdspHp1oVyeFUfm15047kXFD5Cv68OmQPTWmw2KYHuILcjKeyyEFSbG/Vw4Mqjye7lhx+AXvx
KZVNTg9SxsisrcxhLwOYROxrPDnH9BmZg1UwEwibz1qXXRcL39d0JUYHxnPpxdafqV6Pc6MNQlSB
BFQAIM1ZkdjjTkqwarGeCMBZCMK8lSTP02C1qnATXIiJmT9Y0DAp0nUrf25wzYEtwBiPtZ9xHiEg
D7hT1h4uMVgtJ2ut1n17qX3XcC6BdfDHrCqESLlNMJEGbnJIOYm7lFL9HFnCBXqAIMQPUg12SEzP
mkyVB/AMfIHctn5RL3p5UEasfONzlepUN/IHrcJPep00BrbDwNDJaYiQsLgpk62UnpITsHAgbjrh
ZexGdiYY0D4uOFKfutqUuE9pAjuFhzVmLTri1XLdch/Lapel8HZilQm5X5jBEZdzwSxmiy0gaPjS
flgPviLX9kg5lHlyVx/bZ8LgzAs4ztX3RUqKALjvPDvmwcPzeu5btIhfNoWTNoCr7jJ4DUizUELz
KuwejZwBmNXqnpfMSbsUKLZ8lZTwA1Sq2hbqAW/I227MuCCqedlXUJWdtVCXes41lEjR6LLIHMNQ
sOvCIDyKR6qH9K0FpjwLNjTPzIERIqcIaKmXcH9bcUV+Oe0uPvbChx1WZpNX4db2jyt1whdFRsec
8VFGvpiIBWfbkYpHWB/4IO47Pbp0pIaZlPvd323AZbipiymEtgL8uroq0T4/DfXAko5K77g6C/Xg
+lj/Bk5fQHzRXd9ZM3OLTFEFJyHuRjrYzoqUSJAci2q4RHMfxF6JRJLPZBrDYdn+sS8THkE8HXBu
6ILPOwO+wyDBzSQdD/vb6IytE+R6C5lXDg+lQ45Sl+Wst6x4/5pRf75/2bK2Jhg4+KTlqoMemA9/
iFLdkm33z2REi4wZ8Hx84plFpZWTFFQhVjy4bwjua6FYw632jApqx4TFSUcCnw8bbCnlyxiqhvLu
N8yClOWmmWadPSifzm20+kGtEKKrlSrohMcKVOGKC7EcSHE5aCm7hKSo3pU3NR+ZBy1Qugs8b/0k
4Q8aq4OXtgGHys+70MlDOmVPpkktfIW5h+I07Pxyi0+6hyXFFmZNjiGdtUNQoPi5J/N5hL0VwLF/
m1oiGw8oRtGsUdOUeSGcZx3SNrwKp7L28IzbWF/i9K+U+EOcxmvDMAQU+ApaBSDlhwyiPrOQqfHg
BmiVrg8h146HRK5ewbBZqTvXnSY5/OIDoInCQSaZw5BZncyrxv3oe0Rg9G6mZy/V3DMwVeLD68Rn
cs2r8Qbl5ZUjC6FsfoDxfOtUDHi0B02prnN0gBsSbOhAGQQUWCRdiSEpgqCW23tKW12Xk4XoOZsk
e+waByUtL2/Lsj2Fh2wkH0T9XoOVe5ZSBW9pdqT0mTtyVAhZfasG5j6VJoD4YQOrdrs9ThJQIMiX
PQZxnGce+DZGML55vU8uYqMZdGvr4pwii8BXF0EBr9DqvULhuZ68Af3fbHABCLIksh45+MJsYWdR
StYWiirO82s+V1MHPeTj445tWjNNXoZiofBIiMCxoUDkSX9pQCpNot61MN5qQ0xuV09VlcmTB6Ui
FCaL3DkJI9QON0d/R7sTGryqra2jzoQ78bifnYs3IMGqWwAbgXC6MQy9JOz531/hmlwg0HlfyBFj
JnIV5VyFhK7g6U0dVms9B9oFWX/TBTRcuT3NC5HbaGd3lxmz0f3yoJWjqlamSIGYLXb/5IjFHSKs
BXu0H0zh0xQ2CCDBQ2dpmlV0NBfT+yhM/zLEwK+jov4RjQ9QurYm2jVv37xA6efqxwLk1L+PpASH
L77+WYjnOMi1AoEV9w/05Rdj1sYB4egYKbm72hu57LAJpYsCPM8WfZQJuUklUcnQesWR34TGKAAz
CG2VhuzH6CrdL9E0PLo6Ohk9ktwgcN1uEhEipGSgRna91dYhIvl5F8SrDPjKqlsVx1zQSNstzwzQ
1b1Cyt22uNQsHSO5MdA0V7wSnJ9kXXWIbkA4o2BwfowAgaZJsj7UGXLjGcwM99gw4yfk610sGqrS
UK1/xqf6FBPmvQGWfY/xzl16QzTdV9fyHv5Y2+HXfVLE/jLHGwUE6X8ZLpXJa40OwUXpqTpEYYOg
9ULNJLI19Gt8eZGdg8GSjLAua8bboKAz/e5XE3zUHWiuCkguyF2igxLxVtGPTAu2oq2INL+WLJWO
zho2D8JFK2sm5qtpl5ekOZXHgbVRrkzkA59ZRTAKEd9mOy2uH84fzubj1pfErNJ7RmMZSp8nCxUC
HgLtctQElI68Un4KBn+9U0HCUet9A/U0j+MsqJECwKHvamDcceO0YdHc1wp1WN50cCz42FIRNyxp
jdm06X08xJhbujX1J8TVAFsTqzlVpzzqWhIS9KAaPpclnI6WXElqKOp4HrdsOcvZmFdK1xe/ll7T
M9z1a/iMMqGm2GdmScdH3MdZhxon0mGUtRPJQsSeH51EPlvzIUyij9KY/Z61j4wqxqYbABRimKRy
WyzG/4HE2a7XL9QLbiGMtoQX1IcRIL+i/rPAO2gyDPMnxgGzo7rhXBZue/eTW33Xzu51XaWAbDvL
CpW/eSKLCj7lIt+Xy2CmMa2b4jI4lPZKRRgF5YXO5tHeqaUA7wIbdGmH09zDjdpFbmVbJ3XiJMMi
zpvjTdVqG46b3GbVoTrAniWsjpQk9u+qvNsdBXRuyHevRHm+3s3tLl/LqR9YUujRBEdVl7EA1sBu
/w4iRflFIe4pxIGE/2h/Bf8r0ZgpG2n2VTAjr0+gjBaUIMnhpTUuc/rjeyh0P8+lOc2rjdrmpZhF
BIe7T32fkX1o1S3EpkjBGjnz/GSK1xVYxdNDO/UmxhZeV0NoeZ0dePvMZ04Ja1rjcNZmHCQAf4w8
Q2aZWtnrLx43TEqu1p0VE47KVGM3MPq/3l9xEHnOd1ZfQgGbyF1QAxIW//hckJ8Qy2GeWsAK+3n5
fyHWMKkcFMgrLHKQuEl/yMkKYJTDgPCko5mRx/hbFGwxFrHHDwaii3NkC1LRXEsoHAFcabFE3QRv
Yvv9fMF38oz6EQsnEE4ljTaYCDjH5XCIMZvFirU76+0yRLfEEEue3WKDk3TQBvMKI6KuOygRYiV8
QLi8pQ5azrQYOApzacjneKUFmVcilE7OyuZqZ7rMt1QqaxktaT0fMP+DTItUJ2KjyNJfLekQi9Y+
yz8jWvrqZo3edjRLqkkO9h4STGB0okvYFBPTYohCcHojK1GbqwxGwYgInRWLCGgQapmI0uP+fTTU
/xfQIx9fSOA/mapuOQgyvc6/0NbZTq/GvB+ppBsVRGe1oush34jLe3r7XkZwRKPqeBch3xZDebOJ
17Yh1D1D7JqzvEKVG96QVWykR17JBR2AFhBh/Mfcq75DSAgIJTQswXacHNL6AlSg3AtBSFs9dMoU
yCR2ugUC0T9vJQmxjKSpyAoSeEVKJr4GLYCUCv5hFsEameUhTgYknJsDSEkykhlxyNSGtJWfIraO
6NnFx7dEiMiqYXZweS/vu2dWtpyreUeo39Om4hltEL7xHLUHIX/hbb+seqwXYEx+oTYDNVcWkMrp
gsQr/Zg/cthDMVGtSNI5UGaU1QTW4Fwo8LUKD0gkffRePnJWgyPdP/dAtxHHdO2ZfRITrwUdb1F3
0q2EruMZaLee9F8bkZqu5pnOdCxGI0T6TtcA55kUds1geXV4EzycdBe5HyQ9ekq9XkhULi90Qxol
qk6QfUkLjQod198Mo8kSbUjJ5KzBqa1sZFnl3L5O+fEjRSu4lDNtw0J5KX2LCVYFVM/GmW2q7Vhg
mpduIZDrdJWT2ZnfRKLB+GKU1F2kOF6ElTyzprhDRRD/ht59rq0fKOCQrmDVVO0Z82S6pBWg+lt2
D83pWD5+pjutIiGmWrzVXioNbU2fJYod/0wlOAeRqqJSmWQytQzhJED9DUFv11rXBfC7s3zh+rVR
dEdWgamVo2BtbsywHqL2obkT5awVr6s6UxkdIssgpLlfCTm2y8SF3RO18ntmLFBvk2F06kywjmoC
z53YHke0iM9E+BJxL2hhH9ReI6kqF+bfNN/uUwqI49jANrnYKswlv91z+Lw7gf+cs6nJNewtmA3E
kZT0dxP2sD/yB0IeFvS9E0Di6VeralRW+fapYLKbffC7KL/gyDQqKR/EpRwBXyjxlKghkpuVWw8q
TLxyxCRR1Slo62qUVi0CpQw76ATEl3Qx9mCVuEbA0605Vg7XdAKwp9fNqcCSRhuD4K0plaY7Elwq
PlE9pgRZMUrzla07XQpzYBE/BKqNpvv5Ud8yW2ZWk8Y7T+EcHLAglYQmvtVKrw0aBDFcGFrgkbWK
9QNdaw6U8h/XBfKHzCAmKVOXmK3QfQfTc2+XACy42J71qz+iyf8REE17M+DTrSq7t6jIPjUXAzcm
M23uqcHjG7UTuGsennE0IbLWUpZTZ49EgRNZN9+G+P5XWARSZLecQELWGSG725lI3pdj0hAM9a3l
aAg+PR911xidP1u118+6kW30alFwlVvU0qAz/9F0whfhEXeuVtNd7pj6cgK1DNTxlOlx+54NTI9D
6pEw2O3Q1x58Ivag9GC2lQxpggBTHnbE+Z46ih3+cxVKRXMYLSPZ9KSA/s5nrxdGRtRqFC8ebQwh
xQ5z7oD7bhTFjdBXqM6BmecQ9Q3DshogTV/c0oXDpgLkoSrjqyFCd5HZy4YxvBrIgF+lDpeueV/V
A995zPwujnaP3YzPaFddr8kBvHEBw7ePPCXfLe9jlaXxiIOyTOqTpuHhSOYycyvwT5WcfO1gOuTx
omKYaaQG9fXr1ScT+wBPVU+xR+MN0TlVN+FX4NeiJonemPIw66CccRqyoatqIoKOxTBt6k3tjPEl
1wGxLLHS5OB4Trf14pGP/tJF76vESGbHSij2L/0BE8DtquTlqAjzguW5t0Q8M9WRAtCkw5v74UV0
Lx91CSBsjQZJCPvUcPI6pzbmSOzNRk2aulYSYuYmEJ8q4YqvOat0tdgmASzvZO9IPnb2rub5NpOW
OtzJtX5Ag2Sa8fOF7x4IEBJVAhXcSMQX0mAER/tBlWt8I/lkQR9hOBpa+sUB4IWCJH2qDjApi48f
+rteWx2a9yMW50ULFIZ+5utWItV75FZipYcFSBv6ngLq00WrcBl6ySxPgkHKAZ0lJ8/nOkwsK5/I
MYJjGZNKCl9VW9WlPK5XYObh/qzcubXZ2kUumJER543YEQSbKVHbQrv67VZR/JzFKxJvHrKpwuzN
4xTfUT4kBmrLLydHqeJMc7pXQlGp9O/UhIaCDC8YigG2/C6qTTCUgzz5mFFmeHFAqUrkNiS5SfOd
xhxVXT5t2TxhZ7dKfbmTaHWnN9Jokc/4CZI2x10eOIiibxZGQDV/kpbnobAG94WkYN86zh9X0G6W
wijI3wHAF6xuySuuB+lVzdESd0vQLh2XuWUEgebasDrBcZf9JbQkYTFRtkonXNiBWibRddescsbs
zCfGygGwB5l7aUrUDz0KQdcgik3NQ/MxparnPMDA9Ud2PkB0cju7quuqpYw04kV4NpW9qZLsJYmA
ycaY/NI3I+RTzuMtiyXofoN3EZSduTgEm2iNkpQ6AZu38YGyRCy/Jwxfluqvo71N70bhmsGq40oT
M9Fz8v+0B3EpAwqHRZcM7YD5cSdFYRIPLhmjTEx7FpqNFBn7T0HDJP3jkeWYe93ofK2Ad4GVcdWW
nnbCHdRHm0sBcKrslEr8mkUsCnrYZiohEQppwjy+IXUffwdhG7LdZqfYrPDzq1NPoET+dXS3Yaxy
Hit/qAgKHZtlCUu/jT0DRBJ0P/Dhx6B/qmySKO9ThjsrZz8ANKCfYQVJ/yWh20vEU/Vr9LqIES2R
cjOMdR9kQqaW/2SovMty3iLeu02yWRGlhZhAzDEyUw2ipezWoqqKqlRmL0jl3fo6FolX2xW31PuM
0QFgSMYPbECcu+PVPr9bDWVwAjHhLKn/IXXuMxQwPOgGocmcFm5T31yq0/3/i7i9LSyE8l9kCiJd
8pBqsts6UTC63dFu2VR5sRBAsJ12uIEByyjZLQCicHPEXKQrsvIVrKjaiRpaLJyUBvl+RoBFWTKB
Cl1h3oBj8E5GZhTZEGjWN4G/sFlXmh8b/Zm1nByxYpKe7KymUUNmLVEA8CA/n+8PbCAyffVShDWm
pHGgFyuV2waf6Kb472fnqAtmDoNtZbeClCw7Y1Sp9bIlBibb9ZPWlBWzfSTmqBiXuE3T45GKWtei
wbck0nQ5vtGhqoqSCjTWOoQgucBaAbBPqMnv4G2mD1wvBT1bt6kkwpsabrN1mWR698yWpgqKNDnF
ftxFmSmqpbc2Z6Mf/C4+R51o2OiDo/txizQczWGLZ52KP1xJEnyiI2VXSxsBS0cZdydkYO5HVJ/N
jWCJUfKjW+zHVK+F2dfDFOGDS2GoMFBIz5iBAkGo7Wb101q6CjYp6G2YT5yezqjhhV2E3qmBQYDM
jGJL4OrbFthKgkUupLKZFRZqINa0NiDasd2QmZHIR6xV7QF3v2D8dLoRwa/p7WqlxkMYqR3yr5Ma
v17bkenk7Xe3n4l3X3y3djK/+H7ojLsnnefNrIc3F8cEDj4Ncc7wdbm2QZBw+mJQ0etby1SaTn0K
mmUgBjmtcGAkYKCbBHar5yb/dpOcBtFUTqVgyFq9RLsPtQ+VNH6KND18RS8XUaPiN66RLuzlSkzV
vbQQRdnOy3sT5J6N2mqOpeccCmGy5YraVFugt3t0SqjbH+sq6chXFT5g9vB3sRvevrQWnLNZkFNW
Xt5bpCkr1XMflpNuaPGgCxT9fg0B5LDXQsy3OHKvQgJAJNvpyT+DoxRloc5Dxpc9Vj4ScrOLBEgY
iIOJME5o7UMqVJlyD1iImau1TTVg+3qu18sBHsqWXMS9C5bEfJFUbwQrnIHWtZTJMWidHwf64F61
b0juzpr7eTGM6I4+VHfLPkECU4R3mLr5nzkcfBaYsjZDbWWiI132kFnzFxXpUZzEn82/Q5OYSr85
atrAFJay8SstwFBqzqOmHzfT9YMD6BJ7MUTBDH8hwCZk25WkmpiuAoXAbUkxu+39lC+BQhDIQF8z
ghz8zNW4efEI30OhmzMF6g0v6cFT2Wj2uEhnI/Ata+y5+9r6+B5Q3KtAdVNBRWXClxh6ZEaZQGPu
T//TYypANbmBtkaPrWjPkrbCw7TIPKKFPPoqVJS3up0A0L0T85z/fZ8mxl3lQJ3DaBsp5/06Q0hg
LNLBzXwUK5XvgqUihYtC2NHNN/c+vonFmQOsdgoF75J47fO7u4OMWTeVoTXhGYxado2YDy6N/Aq1
9uwV3Noabonqf4Fs2ZSf8ZYjd3Quira0jIe+QF+IpmI533xnxRTADY3C0S3wLrY8PB0LQAtlXBJD
lTsYoMPX0sp5iAyHuXcBUc+DgMKfYy6v5zx5wkLgVUUM4rxa9uOLG8ZRPAEFWIFR2ap9gg89KepK
UIBM9rLckXsqA8PV246PavFDIWcr4rawVOFz1O3IABq81+TX1O1tAsEy8u+u8zdVnQofWww+vBMd
A7M5dKbGPq7V8M1QzrQpoGjm8JOSJJf/iqJkpAGXnIsXW9wnfeHmMJ9zeLFm20WStIv4OyFvs7wM
P+5FxPKltroq3GX62ydahYwfRqxlbinR+6OkRMQvNXJpdxs5lQbvd0y94l8p2TLpn4pSGD0AuqiF
IsYf6Cz9A44bMr4ovEUs01maqSm5MZ24PX+xFQ3qqRG9m/Vx3+jFUt43hbX6n97tv41o1Fbc0Fe4
FWk5zeBKgBnHkagTcToZ0QVzdeN6FP3WtE9/1utFfbMUMHNQjjlMJy1U/IdD+G30FCSvvZRJ3x7e
GsJfkNd49YoPZMV7/n/km7cd7DjaeyrI0HPjKNdaLSkpUdgrig+frn+dwmx+A22SHRV7TkVKT9qe
LOilrKYxrrJImXNjLOuv75fLp/oz3lZYHt7IMXre1/W+TZphwdqe4ngEnF35iTZ40/aURVaZa1w+
FyISfjJRP8IiWlYhpcQ8PFjCseJCaPNJnMbcUIN0RP+msgtgiQy3yMlNqVbR8suH9eO6bc0ymGIy
AA/NMhMEuyFviGB0aiswXtt7WT62y+yE7Ol18XjvZv2d351/SjmX+1MezEzUAOhHjYc/TMKU64eX
TCiKUuVvclNOci49tsjA7lAdZ1vUduJ3c8+eNbZa1m2fQgKjBxAZhtCcueAZpCsf2VxSknUxgUMt
eXNwvufXQ/ltHRHiOA8NpDARCyJRjwdQFDNXXSRsbICjKO5yirpwwVQbOk5jng/IFgaRBDJjyeWU
H6CbY6pkmzeQEDtAyb+WFMYWutufbC8WRHs+yq48uz6Dja+GsCr8mYhNwUw14132W2BfuaaiMnIK
Rs1LwGbhOEJa/uYrHKca+RjUUpHJmPnRIi5Muiyf7GBR2749AdT0nyHVdKki8oRUScnX87GzP9sP
EnvvFcEo89UM+5Sah4WhuwTJqo3y7l2U00nfHhoGEKJwIB47dz4LruZiPPdmQBV3VbZ/Lf1Q2od3
zvcAwflFAF3bLY+OsPIMAYYJWrPztAZlK9i+veeuG6sGBY5v/vRzeNxrdUNbsOPADmmuzS5pEqGl
lGXz1kHMztbkpZ1BOzns3kTxxL0NQ0QyylAG5JZrizcHhV0DeBBDj/F3Aa8MhpaiyA8zFEtyqIIx
YF+xlgOVMPnUVo596purTmAcdCGGvVHB/bq6qpsdeFzQc5oKw/TmqBlADWJLidQK15Dum4M/n/sV
OdkzdBldeIpSYkaUsYsiNGFIJ/XRdIeEkjgHu7yJ/zKqB40Vo3iFu8XtNn1zrpNeFp8wJGB/9dkC
THeHWMDSgA/uppHekw3TvlqbG08f6UWlkJ6UQ6bUgDzVBmBsEQRO9MJeezXavDZW613PQWM9Q605
IaeqwTUVRzrG4Y2Npe3Uc14SROGB9Gjl/fexFB2nqmbt+bmA5Cuu6DhCVuIU2SucB/5yH/2YLLRn
xt0pamL72kt5URw4CUeYSS/x7+O7r3Je9hek+kiII7IwMMv8MwzINlUnOG3LgBhWxTGaR3HzLkdK
OXPAF1acblGApCrbRZwTvNjx+Y9ppDcaKQKY9FusuLgJp4Amz/Fu6NAGiMGkJYdfJupMX3ZqRRLK
krYTRR4cmHcCFJp/eMzkPefuPee0Vh3bXwwcEjN6N8iamFBVRnZESUa5/MQ+J7/6DJTFMObV6CLg
DbKbPH8cEChMZd9e6niQ5jSnYuPiRF2MhzXWtDxQ+8Bge85pEdJGX/HvOf2dnx0MToTdncIuLD7m
UNjCT+BE0kh5BLfiT5LNCe5LBbypmu+JUodKofVc+OShHiT3+qTnxDRZkMRT1Q0Ug6rkA7ID4+Tt
mZ39to/2t9bF22ulIlm6eWNOoS+x6WA/i4J5vbhfoH9TKmZF4rnxphfAeVRCCoSyTPj036+lHkwY
239ZPQpJiJrJvXkTOB1SAuZXnSf5FZtyfMAtysUIpwjYTCIfA+UL5LU03gcrXrOjvojWwwvUMBA7
qqVfTiYCO+nim5dBQprOvsC+CtThFFIhdJBp+y0g+PxcW86mBsz2lFlhg7RKGTvaDsPpCNoJlMan
oHYUrbz1Jg6LDFndH7BUhT16ufxOth3ZZWzMEBsepdJgul6WFPPv/Bi/4sfX1sBRt/VUueY6KvJQ
V41iAT3c+/I2TsubpKtL+FxO2tc56B6GvDXBFbivzUBJLgLp2DeP29vfSa73jH3oLjeUWGJYH4UW
QuA3QYcAAWfFpbDhbz7LFfLAKWnw/HOXlgTAp6J86R8xHPfbUhVLZTnLLGXWwkqi1yQ4fQxUIZHn
GYniNbPh50SbEyY6i/vnIaKHVG5r0gxKm/xYpdmVEfLsnX1lUu4QOjr3TwwlWfPYqQkGmDrEgrZx
sN6kJxao1ehspnVCgt9XXcmoLC9CnnOVcNmQzgHtdtImgNAXk2FZ+G+EayznS07FzPs49+jBpAUf
L25fw9hew3GHjPohSOYiL5FAvguIcLX0hk7ShAE+B8nTNYOlTko8sdDzWeb4H870MyxYsl1m5oLl
3gfLPO49MoE3ZPV+vM9ofScwytCL90SSk+21bYB7RJ4czqesvLYoGCXOu0LhSAP3MsfWHoCV/bxq
I8WsIsVCcRovbrzDNsnCugGv0QxgdDovOkj4rmkrwk+o1JF1Xlu88h/9TP5SUrJFT8ngHpW+dg12
6SWKxUkBmiErjc8JALQk3lXmIT3tnkYWQ4IgVBet8zWgSGYS8GcFBR5S/YKJZFRmdzpLdee5xpng
F7ts+s7Y1CGaoIiXWvrJZlfgc6m8gJs24UylCINwdQqBDxfmI4wq6lVTyD5jlqsDIdD9jGbUu+i4
xx4frO4UdOXga5AA8YhxmBAVDMrhHEiJBJaxgq/TRxQuRzSXBwJE5VgucluCmU8YyCViDK2DxHCF
lNRIczRl2d+TlaRWoEwVpxNMikyOykN/m6ixv1wPjgE59gBIDEYbQb2vpLjL/L5uRfzKgcy2S1wa
UFPuS+m6XVWHrhSGEkmvctow2fCoRsESQy70g6ZrstoVa58Y6kaN5wDxbfsQWVOO3x9QRQpaWIrU
oWG1q+/intfZloZK/GDNyjT0cMr6Sv2uFlPI+v69bNjsablqlFRcr9KqtADVLm8cksAYiN1Eozlb
3cXltgfhAaPDvRfEXKjRo618yKt5EWNC+zPlVqSBi5n3TYstI1wcOz4lWZPAxPAagKVqf4mph5Tx
NLkUTYySbeNeyZtr2YFz8qChh/UPSNSBqN5G8auPTtlU9FgscE1MJwX9xTjeGwKYt14/Nvy7JS5G
UV956Swzni82cc9Pb/Pcwnt385oOFDF0Z2sw0x5PUVEuGMAmYZNftU2ne4O0YD+Q2s+6ecrs9/wJ
LZgVefwy82WD9tGFXfp99BCzDFEHEYRZXBrGP3iKQfBDZBYd3oiPpDyVnT305uFqRfGCck/pH3XU
805birexzXKBGBzR3IYvXHKwfrHQHv8oqjlY6UiZqoWA6lpQgtyZDbNywZrv6Q9vfFReUtTpJFPn
f4+gsF583yetCSvwUlpCP9g3Eb7NhUzZLHjmwqtdDu/WxYsmHdLpUrlhhNN/tCHHNnlP8Py9voc1
omtM2ohZuxhukYDeRP6afBzQG/j/hIAeoNBdyq24kldINi4X95zF99o/qnU/FVH/47SBBglhuyki
m3WX9brdV40jg6oqeaeNWSE0XwYWe1iNokmtY1TaCLiGkrpAGQ5PwCZBsjVg1WJ5fzV/D7oDa93v
fiRXDoxK4/KhuoylJLnSyNiLkv5TMhGMwbw3lALWyfYYNUwpKU4enIY8CWAeXY0Or3hd+Jv2KzLs
ugEjkRD4bh41+aO9M3QCi2y2ZCJHgOx7rTNSWUbGVlY31t2hIDEVQnp1ZEbdVT8vLUdudazkTdTC
zVDkmXhvDCzGht/mMbLa8QkdAvj/i6ojvEfEoYDvPTiF4gJUWMdttIEY8Z7NqB1UTfmeEZVbVDaA
tuwC2rHm/DrAfmZvlFBgBTJQEWSgy/cio3FTddBrb72+V2y9/moxcl1kYVS5QJZBOcu/rbNsbrtm
R8DIp/kp+RtJxoD4md9s09gEG9a72DCU98E6q49+gjjVar3qy9Jo8icod6MmPJ48wxmJqBTb3/jC
3kpO2RxmK6k3+N7JG2GBT2qmMNt3Yaeac2TQeWYHZfmTZXQGqu4VLURtrmS8l1FksiZShY6S8Dbs
aJNsKUrgjjLE6S5jxa1bvfMxnRu10Dnq/sVSDuzmmVfTpMhQBVPJ8llK3qig61esdvAwadUIJi3K
T5B7UOWBC9HaZLlgDH45Td9/p3/1KxJ5zQi0c6AwxKt5LUvpt1FgzvlSUJwhAon2ud3VQqE8lMqA
+yqYEAE7WBv361KPuzKksYDAGGeq3slGeL66eZL2Dbp5TXIC/oXLzAkraSmC+sIcNvjKL1RXCAwA
vgr7ppBYMtssruduQR2+GDZozg9piAH6oJA5OOgy3RYQpxFX++cCLyaNFqKyg6AK77Q1db5yW5Jz
C6u/Y8WEfG/99jF6abNUgbWgBxNfiLkOWEC1X4hfYSGXTgmhjbuoJ0wSPD/JgA9gBBgp0Xy6OGot
azBTgd0cDPB4FHICjHAPSDdDRzhuoNTPAypSiJ/ioHGAgMszJNKlP1fEegJ+y7UDaUzeagrHtaPz
sHPHs3Wjp9Gyxt9kHn2RCT5fYc1xT3k2+my1fiKm57MBN1o7OteZu4iRcTv9IVRA9bs0nB4rHBRS
6v58757ggWpCVlMlv90B1ZrrOz4pcHgtz3HJl/V6C8rhLBbp1RWFmXqX8ttF8Gs+XkzOGinpfWI3
zZdza3r3ZrPqeWrOATWZiGwWuewkfgm21l1MThCKNIWGH+exfDgtgY6LWYTGfDi6WAJKplZ16CYt
8pRcuWZx84Fh4ydzZ/FKJx58CSBl86WQohjhlP7KmeuKlZtw9lTVXiXpbU2GaCC58UleNps7+Q26
733GDsw6sP5o+Mnf9sdrlXMVRU352hcbNk1ePJd8h4eQfmcsnw2C6alKNEtldSCuiVEvAortjI0q
U3e8StgOVvzAkrK2nKqrmBCr2H4jdtG5kQHOv+e0DZ9iOuaasn9nk1QOrcKJHvT21J4FttUkpGCi
tTq1kKRJ3GQ0WMsWXo0XH59Fm6ZX16GWZrYWml8FcyisQ6wKV9SVRmN6uLsM/Q/Xvppd8VkYq+Iq
cRrfLJ7JD3f6e/ZUNX0Q4shTGjHYAT3moVHLrE3kxOdG3ljWgvIqbOl7/jc8PHdw0+FaSdI+hU75
5kBcDTtoUnWh7b6DASCZgpxx82FB5HN+YrbY4ri7kyM9zPKm+zVm6u2TOeSZRUhqLav1o1VoZ0f9
caiz5V66m/naTfARxQmNfclCYkCBsHZLQqWPi48DympYgz26ipSC1TUmJOn+jACezKBNWTRIuoYJ
1Em7Xyox85eAEbHDZT38ckLwOVUyqisZARJTyHtldYfunqnukZyIpsQQrLql4p7wQ1w/v/mTPxGl
tq53oiggeTO8GS7CiMvt25FHrrAafA2W2JDqJb5XamhYrqP77m48pWk9ogd3nRhNrdIWxr5SsrGc
7dXi7+1gpYFZ8XkW9bQ6Mg8KK80JejEXS0yc5ZDS69RD/vnk25gz7+AfE4YLyeNFSHoxuJbelMO6
e4AY4NQ1FItW9bQxtyzG/pMJkQ9jw6B5RHpCMTriZ5TZIbNB/ftCfML/Eo9RleGnWB4tXQX7QgqE
NN+SFmo525EWVulu6//4Ifz9GFY5Hpmd29eUNwyp+k/yl8uEb2SFW7W1Wsgl1XH/a3A8srEassFr
OUSeJHdVX88jwPGIcnHi0dclbvKA1tNwD02ApX7GUcrJX1BP9CbLFtxqC0dCZBCtp7lRdRIayjql
pfVB29Hs6Vk3Enl0+bM3s6mk4NUMzTKBhyZQsWO9Ub5uCseeFk5GOVn94tDa9tHQI/dUjB1HQgzm
0NVnFt3jA32i0IhFMfRDl6QE07hqgCV1A6+JX9E+XV0ZrScqmn6Q5HUiNwbjxHHdo/fYUQsHW7ic
wYTETEQtBpPCyqSoX12D2XGVg4RKI7K1MOa8LuwoaPmKYGAX//8Yl4+hinkYpAY2apVodeySmoZ4
w49sb0F/N40CIbI26LEGn/MSs0ndrmrGb7aWfdn4//1nwV+TWB/BCRaTXDZg9TeV+vDhGAzqJ2wW
vb8vYIZETxYdTAMaD74rtz6yqgVuRQkA3GCFdmUNhU8TYEVcPCMBWq6NM+1vBJjG1FZFPIM3S9qn
1DTAeJsbBeITPjy6iqMzu4vy/posdVykt82AeLJRlAAL+sMZjQY5aztUh09JTLBDU/c7aCy1kU3q
b0QWQF6coeJPkeIWqkS3gdnGUKyAEJLxkU1ho+D8W85r1JaGcxXwpNqc2rMhmTcLJpxcfhri4PDp
GCJIyiwRtT/1yeM6LPy8mgCFAGfYuu0TSf5RSuv0gEosNVhjlJL8gDIzq+PDOY/h4s7Y6qB+n6WG
FJ6pRhbkZ1CRg7HFBHRLiWGPD/EwRYtIa2Qgm10swxWTK3RtEGwwvQRPrGkLRzeS5Pmlmhfrc7yV
dH0hl3RMQIU17yTCnw2t8+EijfMZ58UrWhyzy7Xg3gQBVfQKmNe+dfrdxK9bQSxhKKs35ymkVcDH
jDMtnr+QqkUmPheocmHi4xFBH1SCUnAzzEt3oPZvw7fb9eodLqv8nymXhPUmo0lAF8n0FhhwxuEl
HMGSj9ghvhBIfW71JfcOnC8nJ20XsN+oYukzlw59uhBhQmQs6yt9VPRtdbGhBAcIkwOhaVSu6GvU
hWw+0jmMd0Y+yVJZqIeAFDkSPfyw4HD1n0/mqDkDCvZ5iBl8vX8eqisY7BuGU9/4hC3E7PuPWWU7
tF/1Ab4258aYTx3YzW3VmL9mDoq4DmNPg/7oLHYoRT6AHRLK6WSauOnz35xghzsAgmulvKcnHqxV
/UrmTjOV3qR9xzYFsA4CLHIPZ57DEtaopGBNIrRLSNT8WOiENBVFmf3bwsFAFERSGuhmiG46kEgH
/AJ5+WqUDUnpaobYuR9GSKyQpBDXqHYSiTcFeCwzER/ZJME5OOoixq1FgmjX2IStsEIUPWUdwSAI
GHKhTeZt4gq4vMzxgD6SQyNkQMVKSmRNCkmAHkPEvyYgKF2974LrGZ58A4cB2vyW3+LvrmAFPnjV
3vOzSFwvMQgEQDkdKPWttuzKnWSuj+lLgYWkbJp29j6LDTAKnnZrROThvS4y5qrbE2JujcQ/wAwK
pOuLpZai+3ZXKk3M79MpqMTEcNoMRD3yGcw772xaohYvPtSOK82ZbB4IaRpEqPALaptoGbIt2yLq
A2NmFGyjzTQY+O8v607xiX+ghBfCBELyIsyAGBfWHzMoytmNEjFkFfqciRZ+UFdg5cAyRYnddMW1
o9D3udJU4nRoXc9YjKJ/EaR6paUatjEjCO+eL98d4IC4LyzhNneoRjCvPEvlyyo4Uh/jtOH8BQGh
qUIZRIaX1gvac3E+m3cmk0+RP8UxdwhMy1pKoes/yjoujRM+vTw2LjMWgnTj/g57ktxitJWURz+f
tI+CQwdQ6MKy7IUI4oxyMnk14SEr47dHWLM5Uu4JvVx1Y21XAg/tSd6x+AHlv3NoHz5RbCiny/MV
MyJdRXPOQJP2DirmCYxMBBMBP5O9g+c4XNZ4IHho1TLKREyT8zSVUrO0ohoyg5BuAr/fq/fioLtZ
fq0QJcs3jkukq0KA41FAmPWh2Ndk+vcWa9JFyCoEDH/hWFzmhNpbRQYenXoWZczNyLruFwSBhYWM
dQpMG2eaYzyk5Jz0JbsldTSeHZvWxA+uk+9tj68rMH91zy7JDjg5icv5QQSwz7+ZGY12dz0D0H/P
JmG5x1spBoJuUmtIdFnc2Lv8QQeAFNJaRVro5CRzhyItrJYxwzxWqos9jjFIeF1L7iXkEqpHKoxc
G63Rafb/pdeGqptrYPpXuxbJlFTn7o9/HVegCqIPrUKihsvAlEqBoofu0qf38qXNAx8D7Ov2u5f2
JoWE45cpYDIJuj/fFXSdGi3tRSq9JM1dikF38lxCO1142pPJq/5ybTWlnrf3uyaN9bSpPJLbrrBl
1qe7ejMsprKFcocfj/7beHJL4FDA3yo2fyQNQ6v9zq0k6QTv5kPjgv7fNgAgaxC+ONjOWi6mqqre
qGXdWf2BPuO+DAECfB4lecgN2+N78OQ18M+MKkO5JNcEGE/UYpE+pV+SeeVDhkgkfKnwynEDPDMw
UO6vX1LALSy7PYWYAi8EAR2SSpCfZcBsJZxoVM80ImhqyzCimT6tiyM0F9qpqShiMbWsDBC+ALb2
EBuDvbfaQPl+2mVrF+qwZ6vEdHaXwEcsgL67bgMuWgIqCfjMf2fIdwXTNkS5ca87J8YLSIwWP29F
qyO4bm6BBzD1b9TsFbxz7oEuDaatqFi/HfCqK8mQ3eNybBLm7fTjVQmTK2y3riV4ZOWSswVjIWnS
QRiNInZ5sg6ZpOb7RuuP+M7j5nHRnu7J+bsadtFrxvT3JfW7DC/0CwZk2uCwfwJ7bjNbHzNPE0xM
3lMk/6FJgJdsqbcP+l05O6p/ALM5K+ZID1xOWrowgFcCIbw5ltWR//PL+BFGF6v8GN6qP/jdNn01
UCmHts4mG4sJkmcFHmop1EEbvEChXtBXV6FWtwa1c+R07CblvJAig3ev17TXZHmzWk140tIaHuxD
Yk6Lh6p2zJePezLJou5DxeHLXAatFE25920ESVp4Xpdr9tx9sPtL2R96k0Q4zs1hSX71Q1ZdTDI1
oIqwVCfwRHpjEXzSzhjwC/OO7ENfdyJlJLQQd2RxNuCZJRygSh5ZUyZXliTPbu7vHsj6npGhZXFh
IWD7BgwPPtSroRVgfVNqdy85e2Ojceb++r2SCjuQh0BMpWXlse41j+kviqkX4/A5wHi+u1h8U5xn
tLR6D2Rjw03mJ77LkTm9mOLtgCW1jsEwhCix6j4oBE6IhNlpAadgXTxfHPfyYeZmdImSPiJAJkus
3LUEEh/pnY4n9j8zMyBL4zignnt2sUb/iXmgLlJ7V+f797L4+n5tUC/krdXYnMZ0yivbpk7xtq2o
DDqeUff0nw2xBgOH4Q2glApvO2CxEuRReXpmyMoEimRPacHysTxNlec4Xyt2+Ndl5VBRRvAwRvBA
dnABPkvR6eyKNy7QUqjq/daTy7z5vC8npHxb4KZSseTKOsdky1w4UcV43YmDopzjYYDUEwBFmsg3
89kAdUM8rb9jt5PENtBgriBDitZ5uk5MBIcsSGrRFYT7myrE4cPlF2TxNcgkS5pYLYcGj4QjQN3L
fVUsrpQZv43AgBBK8I76lyhRIGfrfwted9ROFYqxgEpLNfJKNAgShUofd/zhHrYmX81I/D6ISn/H
DAnhD2Na8rDkKhGyPX1x5nGSqEFGHvNsw6i1SScpoWu3pV7pcqhnUZNO6ylSRDD0NYOrESktOgeO
/kXU+0nLuRucKGjl3Df/S4t6HBtzG9Ry61w0z0wwUBmzZB+tBUDfMrkJpzNYlDwX+oCdoMDgINUa
cg6QH8OZoDLx9To9ZgNj2Uc2K6hS/MY3WreQBf0CjnMuH2Vp1htGk8AhUqMfsL6i/rSLX0iu1o4q
tcdQ17RtihNQoKgUo9XMYkd1FseKse1xTukVVJzC1cwh+hLl+aPXtvN+TMR+D7HpSYo7w69l+J7e
RPD7Mth8lOSGzDKDIHdhk7cfqCCVpUJRYQPRhpzCBm0q/dsIkdoTdsUrITztCLwxCNZS5a0h4ZKG
Q7h/2gcro5Z1uAoU56b52iwZroYYHz1QbuwvaB3qGeiCC3prWCXHpUORpQzlj1aEl7zKpNk+IcGV
BqMzkbJ2BDWwVeMI8hqBF1O5zlRKsTzTOTVQEYsfr4r2czmhL+H+Or3AYHAP1g+w7Y32DYNBwkYK
vw8xSKM7S8uYf3BtY99OYSN4P+8JS0mKOTvwPeOy51J1uOtrYJFiNQVaCJwcKIB0bvkZpXD6cZQY
X3TgdMNdMRMtyH+jA5gdYFV5XYrdhok8D0RrDIsukyUrkUtVHpenPsNKlG08sG1zrGj5EuOOeQlI
aJtHu3Eke+3wqMMrsX/h3wNaxPIoB9W6Z8nThZR7wLGqqBJw0osGoAlnDVyut9YQgEXyV0qeA4kK
5pzahyXs2TjLW9745wnFcAtwFZKvPCbD/CC4PMDidOEsKshuBPwW1RrIN8jisxsZtD4dNQT9td9f
t0UF2BKhnqisjojTK8H4NS2MUmE1sh9kNFq2Bv8D72yuV+V6Khh1cxB1p+8S4q6NmavmGnnxTM5k
BQtl6Mm1bXw6kL2rAL9FJHNmWdh4hREcYxjict4FEdy/o+rmuPcJD8Fuya6FR+0YUhm3n07W+Fbo
dO8Rd5XPT/fvixB4GaBWgSx+HoBZIjtSU4mMZANuFLoI6ry2poFf+QaX53oBxZXvl0z8cjS+hhFZ
pFNj84JHMxFE+7HLV5N3JeJ/GUUFGHvGVBs4LOeVsILoriEh45KX82unqk9njwlNUJNMcpUIvHir
YUVuy/o7YvmJf4A4wu3yRKoHf/jjICvBACy/4a6FlQYBZlWV8jQI9QdpCIwYqaUh2ZnPkUTk4cE1
HqKz8aKLxz36TCHfiN1hHkLOwyf9bxf9tNziQHC/aKwj1cTq7kW/hoOhbRB1aqKE83ISYZ9Zu5PG
KixQm+L5fbveFjoAPuHugxZlNnWQujSS7XiwxDYaNq7PSxyQ9XrKcQ2LJU99oBiSNlriPWy8rwZq
krB266/TaiatKBC+fNWIkM6iMbzsIlOihWkd9REXLurWXwm0wFaDFASeVMV5cwl/WmoBZfTnr+t5
C+9aa0uGli9SXcbDkQnlaCm7Z5WepQsMq9xdjgWVY6p8IU3GWx1IasksTu0CMTbhaA3JEXT4oqrU
B5vEcvtQ/ZA0GEmPxee+eYuYDo8n02pV5lLwW75YUfhtIF0RFGUlhPqkCByO9EGapnF+M6vYB15m
q4Lkguj3EMWiG/t8btLQfWOTo/phXjxx4NnmXSTfGORwjl5PUVnqTfEJryuAMquW6Oz3nH5aa+l4
qmHg/Pltd5pSel/VGKruHOwjpuMDfxcW1v5SGblwK/gmPjMjQzJ6rpFRaBjOpwunb2gEAx2tEvgp
v1+s+lR4OYZii29jgEqs/4Ry67ArXc/R4PqdLE8Rdi7M2duw9vABCHoz0qvgTIS5UWul/Lvj5PAQ
IS8/E+sLXYQxKwDOi4Rw0PG6UGU0vqauyOLbsDdAQl6pDDJGQ/Z3lg6DV2AbXH0v8ZZKiAZo1QE3
vH+xnGlkNuxcidxqoEDwVgEHaOeD/JECW2ZbASSKpnoUu/P9mjHCMTf+99vpT7ozyfOo3dc0GR8X
8vEbCKofY9V4JCqFeyTNuMH1hHePBb3f+Id+01zxM5ew637axG7Aw4gqYgIHTl1Br4RujdFlPqXh
veCdkbubpK6X2Vymr+5ik1M2eboRgxfFJZeI7GOYVFyfi6PakGT/rrU8JSejdJVEP6dFSiYxxHh/
Z9PXAwCYkL9aMeGSr331tCFFtTEUPiXaeJEW5mVxX0obg1CFl2diOPwm6teArTL/DT0RRYxJblZw
hdOM9hdaoeD4lR+9wTdyTXAOMx1Gd8tUsDHnYw/BTlu5P5NTnJOKayFULhd/Dd89UyzJRHbO/CkI
5ynBBKxpXHEpaacnUhvtRBQUSvr1FLABqxeiur6iLz5JwG4ox2/BnyQDbaTPPj7wJDqBI5hq9yF3
CXAPLPicrg34ewsa3/4KMq7gVnDoz+4mXcAn5VFgTfA3gBie2P55aKFhS4T5hmJGCYc4acLQ4zLS
F1W94WcU4znlujUFwhULk9fM8CjGQsptrDwGJ+wbrNiiZE0ouNJRQnZ4Ig49kHxEIM7zlS1/2uQ1
5a2Ud8Mg4M4RkivVNJ7xanbD4HL+spP5eOT+gvYUwLtM6ykCJyNjPHkojthAUGmet++4GHPb3Kkf
Afw59nOgvqAQOeBQcSKpTeacq2N25d3F9WMqJrOZ39rXaSoScUsE/6U+67KmeXucxFTvM97WIo+T
6huFBZKiE0oJ5eyWamuCkzKXE3Z3qjkxnCCIBY6alMWRCQalrHBTLy9Zqfi6uTv5SmSfAcFSdBpN
GYh+PTI/XYQoQPHZsiJczWIMXQ7bHp7nj1qoe3nHz8arBznGvyHRjcW9PqbQMFloKq+i/93XvEH2
65PQH+7RUf3E2WPhIjZNixxstbfUOJTo4hcQvp7rAr9qqdbd0pe9YcyFkPRB9Sb8M23P+XE4JdN8
uilu2lS0HXsbpVeJBDAcP5wncqn7BsFSKFJhODSDO7+FQUCEcogfIk91dJ7lfa3Uo5dX9jowpPNr
/rmYedPGTN4CFlk6a4Ve9DcpisuoMvj+DGMcvnTZYN+tqBUgjwH/cVVG2fRus3TeoOfT9WFIm+fu
sZ2Z7FPnD5A3m9RXDZWSH58C4FCe0TqbFz5l2vICbI9XXeJTe51GJ1xBZvjjHXpEgtNkMDYXfYJG
NZEEn1RaS3VKaYEiWVe0dYihu2ZbFuu6qq9byHz0XEKzp5EzRcdlewHH8etGcQfs5Lz/0QfPHSui
iHGJWDFbQnQSXBA7LDQGRM1SXNSliqYfFHtSHpuZoX2FLll7vsP8an+YyXk/oVo2c4xwlAPORkff
YiI+PEuH5RxVKDib7Zkco+jQ0ctfmdk+oM7CiWMmkVd6KcWI6ZULYYETtJU9lRPAqK1RILkiLbln
PVky4yXxHxtUnHQH1Pu+mBPPCwfY6+ObGLYuX8E1KOwzTMgH5CDy1ZlPaIKKBjMUWkPrAhOsTsCo
eXCQ+DjfyOo1MjYXGvdCQsTlFJz90brYaQnkCXkwy9PFAvptHzoc3Ryb9ONU4P70E6Cjp2RWHMkm
/QTT7kRh29xJri2/cAsm425Sg427V4Wp63yqQg6QjWsVXNtlXVbsXlCENGvWehZxImIfdPYk+T1q
HvZeHnF1dIqBEQJQ/De3xiy6FJ4hudmXKoqOd/dsKkytomW6waIbyiRfuncs2TpgIB4T3X0y1cel
a/EFEzdzTUs9iZvlyzFvpcysT1w54YgHZAQFC0Yb2Ookw1XaZ2nkrJDQ9IG3QxgJEUyROZYJJPZ4
HsyNtMHZ6aBapPeoPofw1GYtEozo/hN7z4Mm7WM3wqzgdwMj0ZnOOLOBkjAHKOtwaM68ytomPnaV
0l4M/JoJHvu2rXYdVWnTClkR4o+ILO7/FKtU8HCpQkMKWR9ZlLbNxl0AiAlRRdvkxFOQVlJtMwhh
EbWR/QyCb2v+9J74ojuKT6dL3gIBvrZwO/t7Xr2xUUvlsZbeeNyVDcRsSlzeLbm6BUkNkUU8R8Ov
ki0U0L3qb8IadDQGEN/xunXFqVbxTWD0EIjW2NMIbwhKa8JOTVU2+guWgBFpN1hobDMFH9UwwnPu
goiae8+1PYoeM/3VCXMw6rjgvD9wNdqMQOY/g6lKCGsqhXE0thQRTmpE9Z7M2LZJYkPopYMj4aZQ
HKOfCHEpSr7fkn7QJiD6NWSiraP47rCCf8mb+fifsox92K1IG6eqvkiZEOTiiEQYkZBZcL7h/c2W
aIUCWE23xsikxnmshqn/4iLJQwlmxkx4yyPYuCl2J5WGseHNEE4FB7Mn3qQk4VsFKbYnkmMa+u+/
OQhJbonemhYN/OJApdoj5m+KS48xjFYvtuKTG8dh7X4jvuw/+F7nZYfHnA2Qz0txI9Fvoc+SGMDn
uwaBaA0NEdcDb4aho35qd5sD3aDe5HDCTKlGX2FD7nUXnVPxTPUQ/ZiVzk9HMbOSTKcVXH8S0n44
2IlqZH+MO8ooEeBWQH/m3qNc1TWTeceCEiVUQBJ03dnSlxTAT1EHrcV4/k/OHGFD+y7fmitUzXOq
YUIY1UMFxcIzI+s2uZS8F9CQiYW+V6oYS18lLQeINiWeg7sC118bmNy8cKP6gjcq0u3iMhkBJgBi
S0tQCHZ5qgLfixDJYT97gDsfiIgsqSK0HIFNwAsJJ6O66itmbmIi5n5H0qv0P+vSE59fvYrwDNIR
fPg2iQt/10q2+6gEtUAIjAchlySF8zncReQLsnrIpy0Tdn7gu7/FjRgpPCtm3o7NxsN2txADCF+9
Vm2Vv1QbLXi+1Mhh38V1M557IxFx1TEFZrbwDfZ42urem6wnhya33//XDbxfQvD1koTQLvhBTbfa
W+Ppw0Cpm3TM8vF53WD03E+NFSKchnNHa8dEfP3kndntULJP/uxOwBW2gpr62iPhdxABRFF8VgCH
voaq474LzwFPqBXezT1uezlHGb3ADdS28jVkpQv04xc71uNF6YqgCadGAZEO0dF7xnytyTQfXmDR
dWSiQ1edXP51FodrI7psaDY8J7Fiwflkgi3nO2NBqhmlAFZFqDuHXH/Yb7Y4w1rqWFQYPIhQv1ec
kAh/IVd5Ugky7sTkIWJ7qOyb3HIT9O0UkdOTwZTNykI8jDE/ogMI6r3Mb3KcqHnchQ/Kb0w8e5Jm
RDB7nhEaiypv5FhJR2ZSCclV9sGR7mhHTdKU0s3Rb4i81XvWrx0V6JajxQCmkuXNn5+FBWyzUWKc
xUP43fGn+4JdEjgCUozTdVbn8L6tlk8SB9VrYIGnpeIKXZ7DePR08mwNNhXZU8Dg237ltIurzkxo
KHNZl/HAvOT8ZIQHVqnjzpNj+hH4IxIH+fklZa8p+5cTnK5039s5kkIe/+WnYc9hwNyfwC6JR/GC
7XdLhHp1BJ7uYJlCHyywabvw31HMgVZvWhBG7yEkGCVDjYqJOVOXuMuiODu53k4JbVzW8uC9fTQi
oK2d+QkZsiDd8uyB+vKfGYg2UJENnH6O8XKoSlDTJJ+5oQE+1pASeB227O0VLO/bqRcmAyoMmM7b
HcpYSPUMNajIZ+w5A0VHXiAeJZ1MX5LTX3p1zFF2kYYtBOB9uM0iEJ0WmmeF6pV4yFmGst6FqSHe
x0tdXG15D3GbLly2twoSo/xTDG51KCSwR0g2sKP/o8CSsJtD3JSSZKryKNvZuiLP2sr/uWVbrJXu
rJePsv7J07eGBChCqZWrpse7JyU7wQEqV0PV5QMZEaY9jisJ0eAYZ4QbnW+wMeoYke7Kqf4pyFwV
Z1LFr7cTrn8vaYG8AVcSqKtRKonPb/Q+eLY0jUDPk4N+4qgzZWfHQ3BKx8wrl5uetSC9NanTIPOL
QtPEeYkLmfeRaTiBgTUC5FPlaqPhi4Wpvet1Trywq2yb4ZxKI7ANMBnkDt5Wf09p38Bl/S5Pm0q7
1ntnMTUGagyNaojH/Sf09x6DSAPKqLfaJ5o5feizbSeFFjoMAVCdY0mD8+AK0OSelbyHfM31RrX9
Ldr480rVBJDCkUyNmzXa/DagCnjk3yZjGfR/SFdvO7DE/e9j/y/sstUx8sozZWeFzg+W3VZu0Kxe
yH7RvLxZ4koi8DCKmAvvejYBQgiViPe1t4O176v5CWgBqx0n2dZXz5vNjhOcNfVWFGUW0mnBB1Qh
ifCEzZ+gsQjUmpuDJalz2Odae3akVGlpYIRG4ZnrFqrHttGRTNVSqGNw3M0YPv8ATcYoOdEyjpSv
3tzUu6z4AapaJtRDe/yYHRHrGjrxrXYwCaMh7+BDmR/mVXczQm7Zj0/CBOsHnUfRPkxpzVgm501N
wsdeF9dCXXH7IIGaGLsr00qRfe8YE13LG/etGGw1DO8MNDCd4swiOWDiQt1m/46tU9F/5jqlMamb
KRcboW4GepHroB1I1Td/r17esPQBZnuwwWiGYNI5u7/ICPxZJuYryU/+GBUlxFHkyzwxbL5WW9BI
/We5HZ0tX662m27DvpaHlOOdOdkLkR6ZtOvBDaYWMYYx+zQWE6LFXWiuV1DdW62fOZQGjqFKKvtA
YiXKY9FmoTTtyHlIzxiuKV783W3VV+A5lOGLu8+mizFCBE0tTEbPUqf9dMiL4ftudwoJptfXylN4
NzyVfJNY4oL18G7mSJQQ9s6PN56Ow22YZTOT23oh6PoSlrias6CokLYot4sBjsYi7YDjaVME2JZo
zm8hvrkI1Xbz7gFrpOUkMTzRcj1xC9mXgJv9vdAfxpU1cuoblTTSQDmwb/tCdmWVOHt7ROJDQ0ky
wMXIQDPq0sEHjZ8c1u8Yu16SSNFjwIwTlgPYExE81zVVl+mM7agOfTLUpsuI24AGuj7Dtg+QcKOJ
ivcNimtXxOG/N+KhC03nXvmuNHZETmHY3Ih672CwKvb8RqmQKQWG8wtKlSvEAoFZUmksgd1b3jCI
2p8dMiL+dy/w3Su+U/L4JwxgMejEa+EI7SUAL90wwOj5ity88Qf5u+ouu2C09Z2+2bqp3clhzJMs
6toOYR8KN4iLcS7WKYPTyJrLtfRGgWahdPeTJaUOm2azfvmTakicT1ZpjfUuuKVFhpYcjjc/e8Ej
mXrF9wLgg2Vx7SUxAOCMBZd/aKlz0NemCnatklG8LZuaIawALY8B9Wb5YpDReAy50ocp9TmjA4HC
QvjRoNTPGXvJFCo06o3208YYBDXZg3x5XKvbx1LiGCrTo0ejBkco91g00bHS+1feSWmoyR9ijWwh
8Xsosnn061UeIrGtJfOAbJAeOUAh5FHWeNTtOmlCRU63RfJjUH0LCW9J0Mz9gqCI+01XKKe8gWzT
5ODdVBXBZDfYwx1t59K9QSH7615rErHqIhVhjKOSt1l/Fz1EIbNM/jHAGb41hPE534aPZr7A1k/U
1w1zRfzoGLVnADcmwQ/7d0m9sa5hEWsBYyMbojOfiWOcGlqALC05YhUuoehrxlp2iqq5SEPMFt2y
KEXyywe96G+gYueUimnquk5BRutaMQf7HlI7GAl/gXK2buD6Ti/f6AKZpVVsKZvXSFaagECUdNXi
MqkW/xzcENTrMBE1MJ9PMdl8UNw7+jIa6JVcSBdT8VD1wXVcXO3cw6e+0YbkMdhKqvmLdU84sKIs
vGusU8e9OjsS7B9Kw5/zEjq+triCih4h88p6pCUzutnDDTji2d945e3vBtv7r+x3OIMnunGNUtO/
RxGN3nY1g4xsCJZ9t1d1GhGbjN7xY7VqWJSiCrwrPlqxKqW51pMI8n5r1qKoonW8yE2/hDrAp6yz
pF5Lsx9NAXUxvo4T8ku0mNwTC8HzZjW5+NOCCi2ot0zybZw0Pj2DlGYqywOX0w1QjjZV8x0qbTTn
Kj4mT7Ixk2/MCmNl2BPLKuh5elVxW0g7j8R5n9LWv7/9rAwmONwhslF2TO3ejurPz7wiXTQkTscg
FH+beadrjNFsBXzclrfaSSPIX7TAv5hGuqnh5GRRR0DNtRBecJ8mEI7nNTShkHBNyM8D2C+cajlv
ouvfA4DHANvS9mSzG9i6ilEShgpeLJsb6ouS08QZ7T1PDxmqVbq3pFv0fmWXgcJZzocZUNZnkCsO
BjCjIJZeW0rcuZMDz02GPr5XuyptEDtzOt0kEwKRQRax6GrZ/2xtPcbCW8g9Eg1bhJZlJmSmM+Ue
b1Bs/MLc0PFgfx/pGABjr7rz3JEy6bz5OKX+/4xCD0nDV89PNVqjoveizuYu37xcAGSF/wcjCfxu
TgpMMbv4KF9JmHQdRr9Qad8SpvxIjnDyU2v/DNKnrDyfIsLfWr1uAkxztX3FtIMK98aq2a0r4gFF
4NaYBZPxK7Gz9z65N50/RWl/tBvQm3+hSr56KsQULPjbii+d4bdPI+2zzZgSjPlQjdqrHCN+Sikd
7BnoM/cLWeLBIa9ScLry3VYbR/TFISzqoowIM0iFv92YO23JlGmuaw+nJrev7ZPNbbMam3ejsBSR
JkPPZl7lwE6fXz3Ya4YC4ZoM6t+DrgwCtkAxIJ9Jle2w/7/G80pO5zh2fGBYQGkJMlwxlpG1bYlE
stQLJintaif5Q3aiPuLRNZVphr/9EYVl3wdqboFDiDKDavfI4YC5KDIxOTZSecjXe3RahRMV8BdO
BQ5fWGAWkzHxJgeCq5yOYnbP/Fk1FE7AY5YDxWv2IMlXCWYIiKs9gT+s2tziyPoe/v1D/7LxpJa9
5jZ90nf+TCOpWfq5+th5qFHjxPsKPGCiQV12EAkrevvEcpF36+2XBRz+roHSJWcyxH1xmwnzftwv
su5asA+MPqmcNGxi7yhlFiWErFk+lCoxg6c0kvKY7igAMnXp0IHH00ldCXLLv5G3woCClo37xkoF
bu8QrtUtJK+Ilag+ysr1Fdhh6JI9qG0wlytKuugjN5DjPrJ/rVVYDpoiEHTAPkPvgnwNDwiGRrfP
xUZknH7AN8IO3UVxRGJzaGEVSKbrKUBBY6+YPxd6/5qJ2Nq3/x55BEAVJlcocsw//FzumSCwuIG8
DLN3cLUu428f9RYXLg8h3YNaYY2WwP16qGCYTEdejSkQ9KLSBFcnvXmF9jDy2BTkKRbS2jrHJmFJ
y7EwC4pFSzCHFXEVcyrzfgjQapCZylWH919cC5irEQVSIY700U1OWO/LPbNB2NjnSSLJtDVmGulc
8Puxy+evR0t/BFrQZisErtIlssnbPMspzWTwnDdsehK+mhPWl3CdmQ9a3frvUMtE0VQImOqunVfv
igpVDSw2Z7dpgu98HdB9j41cTLir9eOpTGiYsNe9sPiG9vRSOp/gxSBTdDVZFG8NFcDG6uo3qIao
4odpb+uHXFMnxkufI3axAX8RJ6eF1s3bvWBdWyCP4sNE1cs3wvKCzFWJn3c+UNRLkURsS/xFJZ3i
3tqy+soaQC0MhZHFWbC08IOe3MPWX//C/BqwS9TEVk81+oKJM5M0Roazhe/f9rpzZ2gj5/o7j27z
H2uPte4O/o9NsCSPrM1SP4T5qAAhOw/9GfxZhX3tsrhPAYxQGOeqNKPXmSTBlz/nwP4wg5tPobvf
ddPnZ7W5beNy1Fsx5/XvHMfJKvTfRWXUfB+EO+nL73MFAsACrnH4BLAYhSOga+zSVt2/hFP0BXOY
BaD1ewBV0gkTgmgQ7z89qXolTtGvfnZcoiJc0J9MqIh0OR96+2RGOGaBbK4JAkyCjRCmNc2M+gcz
QRHimmwXdNhxZHFHj9bqwjNfqTY+7EjcrRQCrTpVwyHudNADYUvmziVN8CJDl921FfLTPwwRHZDJ
cQz5/ttMtk5VFbNPZNKhZyi7j7z9tMx/oKb+r5gy2kwjIKoir4rDyMqeXru/28UJY5ZuXrttFHqc
bVf1Eoq7EW3LTo60Cp6Qe8hFpzFu72TXx0ytGu4Fs0jftMoJSgXOR2h1f2HNv70Njqlif+SIxlYi
RhsxRFw58qOSDKTCEnDzA69nTuX57qrTPHGLTJte0VxkwRx7BqS009Lmypq9Mr9gb9xmBjqzxsM6
0KoSOkrwNYC4CCNZfj0lD2gXrJ7JQ5DKNCqihuHJZwyGcXoOPPUrs0r5O9M8sRr65qL8x51BrLqJ
15xJDeJ8CCrXsp5cT/6vSHVKgMjwN3LVAtaEDSTjzi2zH2B9j8z6N0GJmOkIPhL6fxJEr4B2sFsU
7JeM6En2INPikDjED51vUG3FIa32N4u5QdpOZV9K+ijkoqhDeqpAupK5y3miDdLi7E1hgHMK4PfJ
p4RfDjTA1xI1s76M1SqggjxgxAOMOym5Bp/QIly8RCwNloTO5ZBxOkBVmqibl1nKG3YDnR311eZX
6tgY359e56+R2W6moWmV4BgOOJ+TGzti3PvkVL5kolDQE+CsSIPaoIdX0xvqdTgrNqsFZVmXAzvB
ac0UiNhqqSGNPXEAxR+D5tWb6Fxw7b0HSLUfYua5MHq4/RZbHDYp7oy+soYj4VhwalQIFelXCrME
2FLC/31fjztMzJwKukASA1AoMFF0VMYgA62xmhjxvIion/GsQcUDVP3Mgc3LeyRT5sBAFAkRUtqr
G8JDNqevdWpVcPuLsv7HKtgvpTdJ7zAZcSjKiS4iDuyi3Z6zJXg979zy7F8vTUzbDTOdCTvGEHj0
inI34JnIchfpxLvM32BZzFDjo9M/wKinGiuD8Ix+rzUpThl95b/zOIDv6TkajazIdAtrOy7oy6Rz
G6epbL6J8zHbDWTTp5Th9+Mb2p7/x7s2vu49GN3DBCVe1yjK50a9ecFwBBo0a4VFfL/FnWa2PnZJ
v6bBU+AZ1sB9rOvD5qQkC4MDkxDQD9C0b5mVpW5jjDSsjeRDqlucgw7tkZ+rO73iuCVPKCEF2WTS
4PFQFpoFkBIRHiKE0xMA7Bzgr+L238lODw9PpuekOh5uZgqpS0g5ANY3vTZiw4vmlxcw9MP13Ws7
K+w8FenUvGH8TRHuUotia7o0i2V9lAoGQtD2ekMLZjf0ytNB0IRuf5F0OoprP+1KH7k4VC/drV+V
40SBdnYexKQMiu6KMbPt+hhzVmGSmpEX9GPhACF28ugTft/oKhPJMOsWp5oujolmCRt0xX0irVGp
fxwQisPUQenVN6G1Y2h+oIJ+aq7Jgpjb3fQwT2yh9DqCGavk0ssN3LJHaV++AuY/WFCttR74VTJZ
TYONYNzx5HjjQhvG1f5ArBg1UZ0Rd68lkKk+NGqe0mzbSPuiuj6bOtS31nUVJ7z4zDoJVrlgwiF1
VoEgbpGNmUQmrMmymfOiXw+h9Wur1+OerGB5UzQZ8bK0XlDxJKzPhbn8uLE21n4Sa9S/IW9iTqwS
8aXxP2tqeN2skS8BqGVCB4GPloYJ6sc0W7/sWPSHiJwf4m9jozMzG35OlIPwEf+gp279JdcS5oqX
43F0RI61mBWkpVXeXBevgXWSEEOPGTsf/odH/aT0/K9k9UA8A9IAn92GaHwbUId5PIO0hRUJ8NcJ
VprA+UbI2LUharQexsL4QJ8EKmt5k9iUUDqS+8Y9GUHZxMOJnzpjo3JnQ2qu6gd5MztuMNtwDpia
fa50LbAB4z+2QxRQVRGcFr9uzL52Cpl2k+kfcaBtwbxSLNNZ62DJIUamAI+IM8KqTX9ygPYGpxK7
E0/Kjl/tAZFHX6XPcKDSeJ16R5pa35yBoerF6jgbc9vE0yV4KIl8ytFwjKRvVwvb0igL0RYX97Ib
N2vtH4n7XOJ8ME5g/hBAb2sw0eixvbNKZXlfhG0ZFx4tKaegf3j3DcIhC2tF0IHf78QS+bWy/o2/
oVOFq6ao7/P9kQVY5YVzhlQ3Hnqzl9P160ZTzE+sHEdQX9qrq9D5UcsUECl+PX9duyTM+0Ll5Uxs
pBST4k4mX/V+XPi/gDZGF7yqGNAqpUaSh+rXI+SekgswNblboMN56O7ETgOkqGppW6MmHQmzpnOD
L931ubURztsWfcUu6aOxMWUaNZxJlSF1BrleBK+i5o+CQH6nRJXjPtaX6/hn8ocq3p1Q0L1okwG8
KBXdMsILiyLpoyoUYpCaKNE2y1qKQa7nTCVwx9h4vcfWcF5+hLg1+RTHLuLmgOzHvLEkD4fR7yv0
NgpFyRrCxmv7nqBp2cbYF+hNFsY587gyR02Yfts5vLvx3XhoZSwHGBaPd4HUz/V+JqA/UXw6qEDu
US3N+4jD77gI5A7Z8gi95nkv6GV7a44KYZBpyTbht0jFkN9Q8vjlyCxoJDwDaIdwYZluzV7uQg9M
Ul1intvAFBoPIgI+euwJCBhhPi1EUHXTYMIKssrXF8tANcJmTsb/OtXHBT0P268Z7e86ft06M3B0
gUPaRxMV64hXbwHDVL6pzsSLE6DzX8VPEz6sSPMh0yoNHJ41xJs9ujxufeJQJiU0L4T2Cz8+FjMx
6qSVwnDjxRT4343272cs89dzHC8z2YAUaStn9tC4At2klzr/+9YruCnIcM1NF0+P1Ah0EgoYeU2l
wOqhEC2XTmOzYn0O1J/CiuJBJu9edkpgQ3sbtH/3ycrnv+Gh+5fWQhvgKhiFhLIZ19hv750mjlNL
D5MPlirCSrwxrGlVTC6elTRR9g1tc8XAwKhzbFlFbVKSl2ttRekk/il/V7n/KBueXOHnPo7XRAxe
kwZcAHIz5kSzhgZhxlUw0pd0nAq4DeuvkoZlsv2dx4u4ZR2B6OCooDFvwzC1z1E838182LRuqf8F
b44iaO1GIHlCxTgA7YwXIsQgp6P/JAnlh6Uv6/O8rPPF+RGH1zAXEb/zy7YCuO3xg3kPnI8mnpvQ
jAAUZXjOeVm7G5Yel4fLAoYWzhd2aTw0scUnO6GcWZpDpWKToqmxYVfbDcecfzRr3/JFoc0Ugtmy
fKJ1UTvCuVfzAbPcUN6dCAS82rMcCtEOsUuWzjfhLVFpj83OiXNB/cguu9IqpyzLMuUBLLh6SM7l
GvipC+hCKeOpilDR/TxFJt5WZ1rX17LgYdbUhDXBMht0u+5DDWZQLB/APs/mQWkSf7sENmqkoZUb
BOdzGAaVUlP+ZbDbNUAzv36sdDdHAv2UwGWkdX5ZUBJzF5v8s3bwrzQnybfe7SVIio+V2puSVUz3
HURIYQHKy2ABcZc3Tkue+whAJ4ua24N4QuEZMNm7CFt2uDrppXouhF/B248c0ZECHrGLuVqgaOKL
6yp5Hl9stRLqjfwZzyEvHsM5L6rRBYbihspb+nK03BL+A70duqRxOvDt9tCuVplvXGpM0p6Ar01m
V/LZoIuTrW8vbJd/GQR8/6Kw+8k9lIoeTa7YaMGaQL0rfain2AkIgZElcUrjSOp+ZscH4aQHvh44
8ZQJyLG59cXOd8BNQT6y9F1M8OSCyHcEGTWc6Qfou4BswYrraCAOAVRY6wMjCChgA/ZBL2cPfC/H
KfpqiAoTYbOg9RCw11P+IiA6AiPbMpLk/3coBmHrppOeU7n2r9wx1W+UWt9zo0l7s0jc6XUzartH
9rRDnFwBBJL+27+tBbZRhXfMtYnPovMa2mjx+CHnWxecpLY/l2HcCz6h2F9MmIaEQMBcEZCXEjJg
1eg4dQxrBcZ41PpvJzyIeYAQrvB2hegPAosc/ktgP9MR1LSQCyeIstKaQrZuYCV/Kmp5NIRh05vU
WEA20ujUZ82nuuPTMLtgkiqsbmGXFOGe7cNnFCohoWKVHBr3DvouSaIuD0qD2rkXPPDg2AzxlyhY
3sG8dhRX6pkvYUWI6xzl0dqcDetTNUF+Y7mR31pBLANpeAWjJyx3A55Iv6U0LXSTXQ7HTBaAoNCn
pfOquhDabtUSeuF1rrdI4OhgzDW/8GtbOvWiYVxg11ws/vnrFHKAcZLhPEb9dHECl7HYkHhTlAoQ
FgqjGh88km9E3m+S2ykRy1YewnWp9jGLZ0lrCycbXdA9KL6ZDR/j5SFYD2/1PR9LysrhOEjwiGXn
xiXww9Bbzy5J97Krb/XQnhhJNFpdhDAWxqbqUdumHTiznKS/n59wZBJ/bphGziyuwGegv+iyuleO
AUhTEIbujxEfjccu+4IlO7KQLHOp0uyx5LAdsKZ9cvH2LYiIS0X/l6OzbkJhz6VOtwj2uqpPqaQL
euyc3/zED7l4YzXaqw2pIZp5vNwd21aV4j/XDGkKsFV5OkKMkmHA5oa1hpvTZPXvsVaY/oc306vr
DWXlwntJiIbmF7oU+iaNCsXIaHKwQa00/VAstV1S9AkT0gh0tKwjP9TQ4ZKoaLzRksoUWmGe777R
FOnPjKLHLJd2cFP1arTc01AqCqB5S/zQVFKHRXflFeTTUvPJnBwhwmLXVgkDTq/cV9iLknUusGMF
GlRNTtbf85vNtGI2vwB99zbjW9NSxh7bM1ZPbsGhTk+SEy4MEdfA7xTbOplmNydsvZy2H5tzOIC2
oyQZXi8V3oZODrhbkEGy/MYx8cXDu9/lLwJYRsEIE/M3XmPe4L41Nibv6jsHllss5fS5pzPola6J
I+SXN2j6hMaBEsWiilmea5B2tzkos5tLXsrQ8zODuMQBKZSV/jO96iitoZp/jqjW/NIY4Cgo6Cal
/gS8B6GKW0QkdNdqyk54FfRBMWz0zo9TIyRFGQZ+D8gQCz/bkEHB9AjfH53fAogl37xK1IR6ranm
OdvfI5OhdYskNIZugHCOx75ELlFZsWqojfNgIU9JhxWS0oDM0feJbyZ1VoAE4zSf3BZesH4UarDJ
WS22FxQmftOZS+rfL7ZvspbDfNTqQYAYcH40Nb6hRn+Yysi2n+7gQOWYXeyt29ExQKVv3Pr+h9eV
JGQKwn5ecamI4JFmHMRKoe5BuaGoZscxU3cqRNcXS1hvD9SpIFe7/JxOIKGlemX+LGr/LC2+lHtT
PK4Oa7R9BwF3LTQ4lQpGI6F1sE+9FdFiUUOzZoyxk4w6RVU0uXT2I97rJ1Zftx+zo4HIh7k+d5XQ
ee4WJBsoOHDCgyBoM1Nqn5Av2NBIWkXZsmrInaZrgGIwZNDrr40PW8feqohU6Rp1yIvXc3iX25WG
TtPZfH4Oex0w9VAPm/qGegT10LDasD+vyjB1jY/jaXWdq403teqZML60DxtpE2SFG6phpkouoFRO
WlpAOKtyOPm8eO7e9amSsEejVpViSQWNxi8t5Jm2vcql0XN6PJeKly5XQMecvEmCXAwqjBSN9u42
t09taKBkeoCgrBSAzuNeVBC2Kkc7hkifM36OjaoTQ62Q4nGuXS6fxmWfhYZYPMy+e+XLpWOey7iw
GW1JhVaMuxLBVnhBjDJmVTTtjhaZj9nNa68VblsjprEOw2Yny9tb4WEmWDKw7lybMiAjVMorzt4L
RIG9o84BaCWeeSkJGcx8Xz78uhw9j1Zm1+paIKtYIXicrXvHRRQ1fyWZdRFTizeunQoogDgNUV4W
5+J4HJ4ZTvVvlge0iVcwR7sZ0wNjD1+ue/bwUKdnJD1QHL1WObVt0NcWi/CpbbZDkwIj3LdqAXaQ
4hxyGmWjTTuZ59DMohN27ohDR1dtNCboZWZu7ZU5Bu9/4R2r+JOJD5wctSWkhzydTV0MGTJD181l
6G8sJ4I6wrvkYseof348mCAbj4+WsZgmoqnBnEmjD+ojPJ3rEz5caP3v3g3sP0UsgOgK8r19JHtL
NTqkuIWpQ6HgaXD41nZS/orBa3o7YywAo03HrBW7bLtyhk9ZLfY+oqp9ukTsmsugiAPYzewjQ8h/
W3lmd4IU02cCNz4MQBxfhx3PrjAPGXGOOT8O/BU6HmbkBTq/aM5PcKhkX5fQ0kvrlMx6e8ApMpEZ
Ufb60bplbxN27iz3ahYuULac9aB4i+6dnb7Zgobe1LLFvPsIzzpikdfKeY+8Tz4GMvzVSKXVsnbW
GfTw4NnzAVp/k1iWSDGAIjRzFJtv4yU/b+In8vkn9vD106/sfyKq7wjiWh8nsTPQBpjAa4N0oT+M
sdqjoUTzaJA6UjdV/ksTDrpbT2ACObmKaRVDzZI4c9WvJlljJCQLV3nZReF1jdK6SUxSXZYsOmhp
1ospjoPFfrbpTBmyPqlGcp7cKMiCNyKlg2nt5QS0QnCbeyaoJx+NYBk6b1yQbhio8+u9YJAQXenW
OcX2os6bo9KzMRlT7MUp4dJx0Lkh8i9jLkCMOeTzPAyNf3Gm0CoZTzmOzqZmt2fGP8hD7AFegT4p
S4l96ApgOUXOKlB6RyzyuIiAGbfqVhH3lfBXDOer0Zp51iKW0yE+bbfHw//zEbaY98vT5Wwimkfr
X4YSiH8Y12ju1aMw7/D4TTLPdIrFPvChKLlr7DRRJidMVm865xi3D3Yqh03F8xobQL1UgKVb95Np
JyDIJWEZs/6nuhq93U1LmZJq68xNqduCOWW92uWaJy0WUk7nGNLU0A8WXNR+Vmp9WZ9qM0KnkcPe
xB7fLdGGzltjLjpuFuKGG3OOh9I7pYcnZ1Cf897c+6QRePzj0HvvfShYRtO5UVXToBnoTXPQlNFi
M7TUSDGHKmgD5KlvQDRCCmcG8Hm2WMFZRuxEbLijBIKZjAKXXf+kJjVLgs73trdfHvDUSbeB3++a
8eb8CF5drSo/QUafqsRFWfzPVgUBbvCjrNvAaPcH/lsExdQ/ePXry3R9wEI+8AEvEZ1Tgt0HaY+E
msNN6kQPggFo6oCxisguH3JeqnuclLZugRb9yLSJz4XXy7UIE4hjT0jKogccDrTJn6WlCZuLwfG+
8ECPgwdP16Pnq4Ol7BfwfQqa4gYGcE0Xj4hzV9Dupd0HjK4nTTVtT+LA5Mmm3uCLtDtAH0gBcUtZ
vs7ESQQgUoh1QOYnkNgBd/rlW3D6ijMy12OYcxZ+lY9IJHuekwaDxUg6xEGLxrtmI+EkEpwPF93H
4s3I/Ipis3jvv7bNxRQB9oJwWmDWSsCCWY7aatQq5vM09g/LJvNsSTeaoepISVHdTHezHTyVQneN
b9k+WOvSpU5wkzUkvuHR8yn8QY7dSd0VNgaL7jBWWdfBtdklbbUOEyvPsTSSDsHrivjSWaajeD7e
ZZODxqFfQ2uu263KTYV1ZDQpRU1rifeElPDOSKsUw10OLKjjalkNRiNk9EdtSpeeuHq++3FNmmrl
PxcUCm8/DRoy7f9cO/18vKrSOPzbHnIzN+F5hE9q3QpSKUr2YNUDcSBj08JaOR394oUa2vPFWsis
aNmIATp3KdM/OBHobFZ6Q30IGMX/Ll7/aWSv7YnuvMyFf7bzTjK61wVfrfuWRmULBmbNCeMK0moE
USAFNwB7F8dr6NASrF/2++VXeybI5UDnWCcILKBf3wEoTwuirOZyeAu7GhyvQ+J1gBpEWxbIlfU+
fJ2QhQvZJ2RwKu6j8d7Dxg00LUB0zeB095rTO9Bi+oLwcEJ85hnEfBVRdUAWV1c35/KGJxC5uF5I
shBfaaxfNLBZogOldsNb1I7Jda+2FvgCXrdnfjhTeiVIvqBsDbWsxHabiTbqYX0P4BFCK1Bs5kfM
GdtaNBgMiPl6vG8j0M8k5iwpn2AtoaYBc/aDLqbr/+2rt4ZXnNIyNATeQF3wq8iZBqRmnqLhwtLR
dZGHjg4U+/LlttOxzOvIePn0IDqu5oOO6xf00g8wGmtPzVz+/Kl22/mv/k8Aa0jND4IgR1oRbyeM
zBtEHwe+RLNADgH50NzCJ/m+EehwlPI6JQXRJ1vH2O2nLPs4OQB3EUKPda2+LpBdRjmsbZt26pDh
3sC3hHs5fVLhWC1T/CqQsdkvKV4SP0QED/kEYMlRvrhzP0MAcaLMPFmAkyxLXi1kRgKPolsDJaqD
zU+kXYj31UpP8gMdeG97qpDJssIxhgvIfH+fi5c41eV01wVGFrqBuG/d6bosBj/2/zoC1sR0qDWg
K2tVCEaLdlENyR/7mgqTWoSN2SYm5fZllr29AQR6RTKV5o3QwTwGa7hvVfESVcXcjJZnFb44Lsf1
V0esTeYqPepGoKDYlIR5nCRaIKJlojg0zY2tsbzq5EyNLUzmqFaah+OI7e5G211No+VV4NLDAuyV
YuZVceSfckKKbibVPNzVJXPC7jNBoWPYVciqaJVSuGLtYTPV2hEX69x0zhaKN1z0FNLEfn7V0BtY
wbNGsRYj7Wih8muuch4D79cAArfoIa05ifnsMoMjknkdYxo1CIISivITXN439StGkwdqjbVjLacW
g0iIaN+pRVJqMV53Uh4XcxpF1+L8ArS1kgmRBrE+G88jI+szKArnG2LSG/YULZPIvScSBSAoLfw1
oP3BP4dEAm5QvACKGS9gWScN7pNczbcvcdtk/+HXKziTaeR8K2wUaTD6onMFcae8yYf/u2Q+pz8U
Y/0yg2cm8fItWYpPOuLO0l3HOyX87se6nzQvLGd5jwFuNQpf3ldZTmzR9Yua8uXDdmgVSfl9PMDg
wUwNk1cjLF5fdF2/gkhSoLiPZGrvelsHSkhUOUXUDhVlFCIIEJiGYhT/yDb3yD8tzC9ichgeBi0a
HpOsTWRC/b1ZomnYZtaja+QqfawXXUDQxKnj19PKUJu7l9XG9HR/rIOrm0namm4MLR44s33HLJx5
79GnHMxhSA02p13/URmq5YQGrWpNRiu0h76McAZgmhyg18NKIEqJkZerxnLJCVt14Z+IPM0uUXYS
xHZYvZFAvJPNN1P9kOSVQPEOkNAqx/ifOWbmhFrGb/i6953dYATPZ0dvruswV5aZ4iAXE4AX2kYu
yeidmK0Q5QZX1QUlCHTGYWxml1x1bwadTPmMpuGUu/K+SAylxAWBMnqmgdmMHvgPj4KLRaxGQH1t
BBnGTeC4LjbpDVUy0OWwUQ507Sos90GwJ3ALBvOkiyFoBp1S2nU2HqPKGs0SYpDK7Pg2wolqjCwI
18AVcb1oYiwdHOs2M3MzYg+C18URgt50RFhoSwJQ8JVPKu3w5xlwGjhrZYZotgM8gIsJBkn8uUdU
hL2qkXZ0I4IpNzjMBgvw2qEsLLede9wNf+DNgBGphxBXS5e0rV81HFV9RwZF6yHsMZEpoc/JLFx2
Br/BTqjgtbvCUnN/TjiftRBjWqP6wShJt9GvEp6qU0Pitqw+SoxT4XqFoKwf+VSsC7//c/C5kPsO
5/ck4JiZZUOM2aTEFifl18TqaYXZfyE8JWWgJSsl14bdBufpK0Qsax+fSgte9K3TgPnKF9VKIYpD
g7m7fO52z/7i5XecjLC33U00HTBAFdvX3Ac6KMCeBm510juTJ3kfCU0bABPgPE3QJits2QY6vwja
UMzneWggvwexUYzrIZpNmOA9dQBebtpGmbGRLH8Jp9nUsmY5ynRT0a+Lp+1r5Zbcoyh0QIb5ewKe
Sfl0BWIP67vdwet43R9Pt3KKmN7B+56tQcz11sacTRS7LgJWmGasMgo5ZdMgEBiQ/CkvWTRCgXQG
fVl4+ZsTmulT9t6nqpu/7scvqrNKQdZk5rY89e77BhJstugOf2LagVKiPOvaUVzyHjOCe1phI0Kb
OU9FcrWNxYldr8cTwxE/EYoaYgEgtRncpXozRnXCBfTh6wzOAilcwSQ+8/xErktJK1Arizm1J0qj
x8JyBh62xgGChwe3e7KAOCNgMv9XmrC+np8Vp0f5ywQDqsmd2uFusMeM+/IXcXrF1kzriv0Q4fGR
DAKGUdjsKZM4Jxl7UwDNmdcoqM/fDlyIPFoL85WOLfxIURV9dZt/GNLLr0uOABdKPSiMX/o/Ho60
MJQpuFb5nX+aMWElhidRg60S+ul/hMJGgKIwyrPf+z80a+Na4JFK2a6ldvdBRr51Ia1TLIRuKNZs
IITktxzgQHR3i+klOeEmSc/L8fQoUwOS7hBg2sFiTtBAPNQOxy4rzFpyLmvbZuHnOeU3op0C6fdJ
MPoelxagXz7S6VwKAza12WEItvcbRtSbtoNmWLUIHN6MvxFx8ybktdKTsRqNK+fBHUvmg04Ad14P
/Gz/mzXsLsijaOkN5/lQbrxiMNvwtajN1089g3hFp2ayrvHC0zLILjVU6ZpWS7oGUulEE3W8f0oL
dhyGh0xeqRzZcVh2CIxwAry86VF9CP+I41tnJhQGTuWZg+AFByIdkfHtli2+14vtjbVb/pxCit05
xnAbT+1YGA8mYEC9HB5dT/mvJkMivKbmjeZhhT9i91yKpknMRfHlKg3agy58pD55J0cCBHZcZJ5d
N0KO3CHdsNUJuqrepIwvDySKc585Fs3m+5YsH2n9wtZdFjYc58fDioAgDal2uOyPz++xwVtxS4F+
PKCAoqR6gdK9TtuJqYKHLA9jMi5UgXeQ7BmJ2rvX7lBUOMWJo2Z/r9+BW8m8UJQ9NESMYl9x+7Tf
t6bpixUZISyC1wNRSzl6jGT/4YTD4hDijGAYS5/fXESuwSpzSr0/zleqbf2B76QYxseiU0DAKO9B
kSyrqsfUEF/bRFru0BojprbK6BXpzI9ew1oS9LgNmR1xyJPPHmhbCUmtCpds9uIWP9o39c1nx/Dp
9ze6wd9cPerNkGFHzzAfJGpiP+TjlgMlct5DtkqIbUwb45du0HGdmaX1GcFjYysEkbRS7WEFcXId
/p1NjhC0ZDST63HCWjZ8OFUft3OK4VIQdvIzz7p9/olXdtdmWy0PYmgpRq0hmqfo6wDILSvY1SGO
bqxc06H/K8QFkHKM9RbJ02kZwRHOghMq44StlvJxS3cDpWt8tLnoS89m/Xgm1KrBKGxYmHjkvNQq
fdfF8jlEPG54x9NnL01NKFzaBonaEs9lsRui8yMkvASswC0vxNe6fLk4Vwo1RnRV6YBg4TkHce13
phaQOTYLh6zQNIFKBkxvLKTvvOeZOGmt/GEo4MeB2dfq5S7oUr4a6YH42jgrOL9J3SLDLuBF5lZg
h1PcDTPuWIWfxqAC2aLq1e2NuIOSJ3qe6G7JBNbiT8LTRtMkHCRBlu4QGoWwNlbffaTUex+Ho+Oa
h79tvGRzv/rWHMTZtWYY6cQ45ke4PfXTXgAnuOB9Dh0siMEPjXX3OP+ela5IRbhU4IHgzd2n9coi
2uM2VwkcvJ5JqzMJq4t9Z0a7KQqqsHv5kkI8aq25VY2x8t2QMZkIzl4Kwa9a29oEqyE54vKfbAo5
o9IRstedrEj6jTBNenyM8W+ji+lHpgPO7j3Auqgv3/aDcmjLaC1SdkEXNHC1vFpAKpJP2lLuwmTI
i3DIusuhog7iulj0Ku31fqvpH9DcJY7HGqJ7uEYvbzgCCmTtrk94P25JKs7f59gJUxYudU84S8hw
oyXBRZYGM5qQt5tBvs1fjdnxRqCe9ygeC8e/X3tiKGSggt6WFWw13ZhbCw/8xR4RQXbB5yHzhYkJ
ptZ2KSCPz+N4QqOlp7Jjo+JqgsOH/ibSqa50InkQdbq0t5yr6g3ZTlAubNM0+y7/VjiYbd0OwiKx
6hOq8W0gcnWTt5cv5KKkr+Wd5/l/3xYbEyooNeS94z2kh71PswK4fE3FJaUQV4W3DBoEzT6bGHWk
UmPGSOZfABgr/RukOcTthmd/96c4/CZeR8Ce9LgsfyZGhMg9N9EyHVp0jMyXEHPv1mCoPtJP9bzK
KFw3viZIFBhTjHl7Gt5xKRBlfik+8PATS8PevhBg8kWHBC4o8ae0mYtpBS/DkfUXVZdYqxsXNpgA
4tCA/vDy4Lun2crXPMjZBC5/B05yNuN0RPlHES52j8MloWpu1PIwJrSaCTSmw+U9TV5da6JjTydL
qpvKQmkvo3uAxwXetFdB4qzWzUx5NPLJ/bWteLavZs5orx2y3U8DiBEWROGeKymVZzcFCS0KVgJQ
b0vDhF/xC+EhMGRV1i0UKjWdOLhdHHfoCaH/0ncIhW0Gr7V334TQ9waEz9vKZlgx6tQ3o/QMrf+q
R88Y0YOasaOREt36R7CG9QuA8W8SCp2btnLolvT8vTOgSf/ZxNFBVVTMTVitH12ex9PdLEGB/7qO
P8UVFdoUEzvwLdreq6M+wsI4vJYSXL3k1bEp8JvUWHy0W625W6B4eETxaLsPtXhJNZsr4lVSZSfX
n4T51kJBurfmn6TLxkC6Knhg/cWv2OkqpZF8/gW7DqM3lqd51pvXm4nS4yP/xYePGCKffZWH3Udk
fjZn7s1Fg9PMi18jafl5VuZMen6JMffDti3ImQAeLjzuEnO69pll6DDjAzrABabrSduVpyJZsGkS
LV5OA+E8m3ayDTwZVOh8ZTTVGPVlw8ObftHqHmr3SD3Vu1CmVyYfyiLPJ0QT3iyKjnZAUqPMfl7v
7cehpmXFscDb1/H58ERM5/3mq5a4Brnv4q5Z13uUcHD5MLeiRHu7x21dBY2mGwIxRYbgF+75USZ8
VVZsGtvCdFkyGZXP38uD9BFuGoccMf8LzeANlwc4SzpbhFMKc0iQcIqqDeqKGdWRxX4oa4fMOYig
hlPOQdVX3bSfettm9dHfzGqLkQ4SKmvWno18jFB+i8mgPDT4zGo8hTiSgeu7QChyFZR3orcYAgUh
MrwSVeejLgXG3Huj7Ivx8VQW1ih0vrbdZ0ZCE7c/Q9NwXaj3RPbs9YMB/x7t/cJDYYCOGwbICPn3
QhJ/o0G5Xu7pH2v7VYPKdh8Z7c/4EK1r3oacHyJhNvfOMOJKB3wWkD9Ggqh78J96X4kO/MV6X3Oh
iJPH7wlYV+1hrwPG4UyZ82ELLhQhdec4OUqyL65I9QX7AczSoA0QU60gXhJ1wFLnumdVcsGxA05J
CrcmzeZuhvVmf6sbqZXUcS1fFX2te5kOkIJ/xcwNSm4+D1GGuKxOzwPrAg493781wQ1aHG0PkG+Y
xm7BOC1UJy7YkIpOdnE2zsLNxDzYMv+kK80rmE7fgvfplkhFhSu1HoK88xXQrMsfgtSIY3uzTjok
OXDxcLS03SKcWqxg5IPwEasHoyaZY1FQY21EUxNjOFN/0vGm+Lu+Ve+YKtKS7tR/1vamfkc59a/d
Zx87xCQOOpZOGiyVT4YL7sChX/rhsG3OlIwbTvXYGinM37j0trLW0EqOuzYRDtRQhBhdx7ixvD/E
zYiERmGvNcAmqOTCWNe0UQgs741yGHqPf9XBqinxnZ/M5E0r9xgmNezp3jrj158U62s0SxvEltzs
2lf5rK68PVp4P3nqyApAwNiTIMWOPkdw16UUJBHwb9QQNZ42AUXmLLSj4hxH54odj6djp+nHZDml
GVeTFl5a4ilV/L2hoGOnBwuPBax/Ke7gnwLlixWvPrfnDt2JIGPIkbrd+qALpbCQ+RZbP0hENE0p
Etc89B6VUrzobvSRfdI+a3rwHJ1y3b1YJZQ5+JUtqPqugAwM9Za/YwRebeOiEBO7LQwpi3hSrUa/
MGQJYrEAeeAhVznVbicefvKUa3+tok/KmgUScBTVzzw47Vk7xdurEwDFAAnh3yi2iPMcsO37Em6k
sGaHi230LAsikKO0am4490i2ehAirGwOn+6O9dwWW+WevY5GBiqk11pgC7wUoY5TGhp2e7PEc4O6
OW2cVeDKOg+euxAIvQbxo+Rr1orAauLulzuGU5RakVZO4aZnuOEDlqEAajMiB1xg2QffHI9N8cNH
ePAumE4HSnv72f+QHgGrQ8i4AddLk61gUrIxJ8uWxcGBG6PO0c1fd0f3fm5ztZbhtTARE8Q297Cr
S7jNZQQqytgrO4xelAlfGWWr5u39p9THbUwvNFS1xPqCIA557MyrTF615JoyU/FPVlK6r65Fv5Nh
/TJQpuaaVA8dVTtM10k8Oa4b1c0eIsttf69SQBPbrG8HdTOZ6I4wcX1eQdsW64SkWgO7GpKsHm4k
H4bD2oO2j/qOfaFWDjBy2yym/ORjs1PdcHg7Bii1P/d+ggO3qQJVE9zmi0dcNvC8NXnwcr+7wUjO
1u6/HhSpNfUUocO6dJEHa1MhflAt9jwPBii3xmacYS0QIc5zU+EeB2t5+lzDs7PSSXxkKE+UHowW
CzSVqjPkbCft+nW2jQHUfyRh4tiH7Hn28MeCG9RZJ3vGxhKQkB3s2YoEMIlBmxUbd96szqf26yYH
IcYJtdd+Ch8Ay4jEsWgPoDQ/rnXjMUpCaiKnngi+slDJjjM4sHrcueGap+JuZQf9OlqRsx8bswVY
y3BfDFnhlFuebCHscfysGZvVe/WBo85lVRUCahd604PMm54YDTULj0wC0xuMohSykBWTUP7LtDaH
YhvhNFge8acFYQE0boWSCABuMvudl9wUdaUGB/Fe7FhdmLQ3ONZEWrnQXXf2u7osCPpPI/Wa2/4g
Xaf9PurvVUJYbtfNFHYgaWOHYqAyoEOCeHCTW3ow11oBnB96H00w2sm9/i/3yHDopq4kVWJxk+7A
PR7ZH7TVlMzenQN5BlkLMVE7EDFjHYrQn2RwrYfdnznTlDwhuLDvDRQXe+QmrxBJSGSp++LSFmZc
k07DKSMMLPTNSAMQHWyfWWMQCdZxhekMO4H5E1wNK/O6PSmv6McRvgnPlRMDYUWuM/ESVjl/PklS
xyLWUIL12R7X3xnEAn12Khl+PqUChQV286nbWZhZZ3EGZRWGWbK1P0lTQcINx4v+Us2FV7+gmfoV
IHlEUplKPAqD7+LJNtyR7ZrRT59XzxkuMMKNYqAR3rWheOXaBkGptPQHKu0UwcBLpqLpK1X8SAVJ
2uviEQlErmsjSShwM2aAvZUxgSgbUaRLqyZrRu7vbFR23aBnQTDuZypjdelct25zYGMU/GQkeFYX
yCpuFuI1M0P20iKLQjM63L/dsDpEM2OyWnwc/gAaWYwpzmloeUY4YQhqbotCnUylZmkbI+obenyf
p/g/+/C8+J35zkeFLsoqK1rM1ey3gIWWUzMFG8LBnNxfmZU2sADw2PyAPz0WKw2XwnviGZzspjyz
e6PM+dyPFjiIhBzPG48iowIpmIMqwZSo2Y+py2nc8UQAV7whx40VYVpOQAM9RtpcZUzx0Oq5YWQW
VxTIbfwrTqFfRnCcl3mDyfLc/p07JJo+8zRftoYfS8oLntH2NP/EtAk30piUGjdFD6mAS6BOqO53
C+RTRLeA+ZOrl1W4Zy67PhXoDawF9IQCfJEaoFCoawCXEzmzs/bgKIUDzDIjT7SpKReXgoTryAzJ
R6qJa2mEGBsIXB7C+/ROKh88DCHhvSatZJroGpjPPihofMaLlkP15/LGSuFdlzekB7oErzjH3NrC
uzvKZJ7gzCGC44a3wV9uxUQUncXy4LJTmzHEDUibcZ3Kmb+kMcixyUSRRtp1x8ZDbraTGWaJRraT
VNDw84rA4um1UDnbcnSabQkNVBgRXVCCNc+SB8tU+D9wfkGYBAQq8Q5wynyRTvgiPOZwiktFcbeB
qo3iRxMiQIhzDKIzUEyC1jHV9CuW9YnaC46PVXxI6dZD8F8VaPQw53LcKWCqnHUgT6tIodAbymA7
bEc6M8Eq+Uyi5oTl3bREe7/JjeCRK/hjkJ0cTCy8dfpJIxcun4E1+evU6YW69K/TypysRnQWHGEJ
gOwujo7NdyyOLdcWY1oYsZprY+HRWU2MefvG1XwRN6E8xXR+iLPDEVV3MxqjFOxqe/ezd1/yn9TV
IywePquhGlHUTh2rgyfLNQpY3BwvyArwa3UHLe+5DUDfvqvBbj2E5r2pGy+Lihv0aV7kkXl59x+H
Fl0KmIZFLbFvvdHBkgWURdjwzjWiO5bkqgbVNKJhSQ9J2/tAl4aX6KF+ceCYiYJelaBlEXdGhalH
0l9g4whb/Vh5m/vo1FJlqhHGRhXNuFiQw+vT5nykRGTkmWU6xejIUzorhkllaQJrymoXamSaQaqC
eJiNTRpQwdvbgVuELZ9bT8Zz7SDz3Y0/cjk2XH/Qn1pOt+fhzuWUMGOsBt21KUQGvOxpU5UwIVs+
zlVmzatUY9GIlM1nQmk4Jw/1gRttopqbtcwZNE6fV6FBnqQtDqqYKH1aF+EZmZJ+tNiXtc9KQdDj
NFYekX4kNN8Vhd0Kbrzz1rVpVZWqBuwyZUN0r71U9TvluZXHPum0kxtKzDIXZWc5Vhiff9ZeILdw
UrKagd6FJEiO8M3bVYojk4X651S4FDTHYLpKBvOSIv7YAE2w7v4HTkWvwbC8DwkVDX//uRfUi6SO
V4NRmJL0OaB/E9h5VIBtkN076xEeutCexntEu3KcgQKR+BBmRCcx/9DMTpb0trFDDA5UyFSD93oT
+e0odK8Y5x83ntfFzarLJtQx4yqCJxO6F4mlzr1FhDInwDtoLPaISWL6UvCQEDvXV5AG3CWRe0oY
Cut7NPN6zOQ9xU8XuFEU9yuzXxHSAwe2Kl+LyoSGf3G5slNQBMdfjvwN3C6ZGxr3Va6CCdZvyBJp
qebdg5oNdGAv01sb0lny1uPu7XgoFZklBN/tCAUVVba951AC+YBR9I8pD59IEO1fLYxgAP/w976j
HKEo8sKICDzZECO0pjaZlt+M4SBbpHq0EYwCY0feXm0Dkpg1DhImpuEhh4Uq2UeYwAKBSsBILcRo
zoNL1I7GtGWUv+aO3Pe9j8JDpRlHm9nPJkGxHrQHdgi83lcf1kS29ZjHU8WU+X4YCzvoEST96mTE
rlEuAkntR/4guQ4um2mJENptTkfry0pRD6Yys7phuIU0dadFMkY6z27VEq0lBZ21kzzh25IbuTAq
lCiZ3e+QTkiZ+EnFre5jhEiq4lV2RkPeufQ5wtUafv4XYDNQPy/yn8ALRX6YSDyBGZpw2dEhxXSq
rYllV//JyUtT71OskUaruOKyFRHvbjuoOkZeywBhS7CA8s6iGmayBJgXiGjQ4kSHq+ooZS7P2cxE
IiSYHliQaaEid7NVDjcCnW6Cbt//H17hA0EZGH5vkq/k+8Viu7tt/yBSqkbbzxIP1RZCp/ZEU1dg
94I4CTJI7txQxRgUOuukEdPZygOkc1UYQ04r7+PyK1XclMyKsXfxn6DFdaXX6qj0+NkCLe5qjX9p
EWPRIpBPgPPZ9Us5dhHyCx8t/Sv1dUH2iN4JYPxfQ8grf6T8nuKiXpap+9LplJu0geS+0yMOXngn
9+MWj9ZUINj/6tTZOovxBQQMI4f1UH+wwNMzisxyRmLI3WmVCuHxt9aLdTmgitz9pNZd8vncPqxF
HWkC6fA838kXs7B0xeeXf284pLOmtwA2XjLzUSyqUmDIvwo8+OPuuCgwM+SyLZtneQL2RYg3skRn
Kv4CQ1HbwfZIX3uLfl5BnsHFG9aVoZO74+Rp9z1NIAYtlgO28GR6ojOmqCz8/10/v5uZSJ+4EaJC
rXCOZyweFjsn8UfpHozx/JR99rNlWU6ZrfLs+uEThSSYKbKp1HF2SGFC4QNcNkmE+01P9m27Wkj5
ygNRVi5O1tmNJ4e94eflqky+QLtsstLEPkXz6Ej4WdJQq1pPU779rGQc2NfK7LSzDwPuE1FqdHL0
uBTvhbBNKCMg/XxG5vp19JsYaGGAbvgRcH42En2ye8iWpm7Fm3FdM07xv6l2T3zNeOEmNNQ6jNha
2L2DNDi02IEo1FX96FiwYYPYU/cYWeClu57GYiInPbg9F4sQ0N6Y/8j7Gapcv6RHV9h1e1sJ4omp
+004Mnl2QZD4Hs/r4PsHyNVwQ5nvrHDR8WEOnHXgAfXrcn1FBParIQG1/sNSvR9qY9zg8kZ5tzyj
4V7QgUoJLBks9MqpKH4tQApPpmjQBi/BgB1hfzJBl+4sV4cV5C0WxwDnNlWthqrUgaA5p7bdXo5f
7rnPBa40NvH9zuFEKe06qH93GoPWEK26VptbXKceBf+cHcaukLeE15wV/GWyX6+JuPxwBvb3smCx
bR3CTOKtrphI1D3IrCDkGay9hdQyfxtmn7Whit+EG7R/U1wUr0VKo0lrfm7t6oRaOvLzdAt6p2TO
ImIgtaT8SdByxgGrz2easYHkGtg5Plg4FKU9XL8iV126qKniFDD/2clWrKOE2y0QVFo2/Vk6LvNe
WYw8tDC16YlGqpr3qzvd+p2riXjA6DqJWOjKuFfTPD27i1hxV9edbvHGPRReG/iRdHV/8U00ULek
/CoGVsASoItdsyzihadAiBBWo4l/fyhtZ2x6OWneo/6KimuYm4ypHi0W/Qk8g7zo/qVHTWJjLOlb
JrzTgq2nnuoQpYN600Wf3cnmW9GP1JeXHps2fTbkTsZXGEZiKsetRMQjTe1U/kogAIq+SwMTOZPL
WoiY6KG6ziFoqbEoseqnP69sMfrqkukhAUtFrqtaIxsdKhT7FO6PFbtJNGj+q+NrVH2i7QkdbSoA
Vlc1yi4sjb108inMgmeIAoo4vEHKmb+2Nr3HqqcqXND/5q+IcGALHSE06cjZMmblFnhqQqeCol82
AY4o1iaYwftaYL+plQtPVwhOjQ1gzG7JpdmE+j2VFv5LIhxj7IrpGXddhIW4foqfKmAnr+jFB6Zm
0csN8cYI6im0uC4jHtg0dfXIbhflS2RVGN02I5YIXXyWTuIyMXODCrOzsXPp4FIYJQTolQ0hxaNb
4BBRfyu4pE30r7dYEqI0LykybvNO/7NRm6Ai6gSITTZFy+7/vRWNXW/LGSZqz7wWdk+wAYtYjTD5
HHgH9qCsVkXORVw1i7QHTq61PD6LNjlWvRkUv7OxsoU1U945bah/g/vIjT14YPYrHVc7J6FVO3nj
ztM+A76lZvU+/Yr8x5p+ebxCHlRTEZfczlz6hpJZX3WYrcV0wYCdbtehATfSYUqDhXGEsRd6pnFK
Jw6T8e8XbT5got3RTEdoRDV3RSfVm6JcCxyyEecP03xCxEDftzpH+U3XdJKVSPhJhtUIH+xzetfu
ndpNuB0D4BW2Kc7zFU8tjKo52PV4f/OYl/ApIIdINAmSOxhUrxMiaeO7TbWBCqscJqfSXiK+swSv
7QMR7A/oMWW0Z9XdV6HBHUTjUylyMw2KcU5onmWxIAMz6xH8thExzXqCnO9rycXjkJoY2bedIDs9
/7vyGb0izXetgrD1hZIoWiN/DeZkscJFNRDMeQZrTxilYE+7gApkDrEfx/ODklm3mrBwi+wCtGwQ
FCQH9V/f+WQlEtU1ohr1Ty10X1s1NX7m8aCkJ06QHm4q4mQUI940yB2CQr/h50//vMyl8AFxF/2k
OqGOAb6lE5xBMnrY6xa4tIWJbeOvG5wwespsoCIgpEEzrvQWlUObjcNaXxUW4NTv5XQRUHnNfKUZ
Nazzcw0CuUzs7GuYtWtGNFUKqQY46+E73SC2wN/T46dgNlOxN00iGDabvoNQ9REgLCMA4GJDxEeA
SoqcmAl1HBKlsNKhwHcSwHjXYuJRCmCE8i6X18xeDf+pyp/k3X38E8zqPMGoxWkgvdZ2KW7d8pw8
WKyvCMVu0BlMTHQoxYMKCRTrmA2XVs0MIYDvgQ/kr85qK0uq+gfP/aJDg0uTgbo4L2bFq63+q+mU
rrfTMAs1WiQmqks6Zz9HGOFGWsBCAbmOwLVxVBWASf1Iu7RNcJjxUmFily2oyh7W1hl68JIuh5zj
Do7LbWsxexaD228IdWDxBe9bXc3W3VBZ7WOO3BArE9D1sa7UDbvt7xRB64X+sDoKfI6PChcKOp4H
orD8BWMi07rlTEbbYdIjR9lzRJ35xeg54juISHnl2XVgnIosU2Kgy+z36lEw5DjT4nqMNch1joXe
+Fv4vRwBZvrialc1gf/K3hC06BZRTTh2tInBtGlbv486jSTSTdk0z2oGKxRJ+x2x20mwSVRbOrjq
tMNVx7u6vgevODECwmrTG7lUc7H1F8O7H+COR/B3LFNc55WckIdlMri9ZfTeATPB7idl1Gy3cF6M
9mmjUAUUuxj/ZKFPe667/dnietHTBhFj0uAInf9eYCoNRfulo7oiQzpSwX87I9wb/VPKWneQnDA2
XBkYkFRA/iqQLKx2Ko2Iop1dn0Glo/rSktTo2tAZmY3eMTt6xdObLe7fjG7weMRHPLaO+WfzDUZr
ssWSDIRKZmV95H29nkXsiDxGm0g/GY2ngb1rEgsaubJerh40Q1irmko9OVOV4JL980BIZyAZLFh6
YvQAOxRjvwffsEZIgM3/ax/Wb7zKfqB2ghDe9O6wFxWpkOjP8tlOfem6iQ15p6A52YSxtRiZxx5t
L+qeYhHkE8cyoo8YuRZGL9ZC8Ym52Uai1rHu84JplJ5oXye4Gxw/zeQD809Ru1ToJF2nMcX8hhte
7ssPfkDvZlBWq7MmuggAKS+TEgSjIX+AWo4CZvNJrBK4dXhDXHhPlM0qQG0MRKV6ynXsZ7gvKaOa
Nl94uWaokZbwmJ0gZYo5nJfhgdY2IeiDW9U5D+gohHrTI+HG59xraGqjDczCUcELWHw6iePUdb54
ylHKOTI4Yet0vMKvCbjnFV6lBAL5QelEabKhNxQmDPSZErnZgu+7DAmFTYoH3RkSDbjm0BshIbDQ
b/VjxJE+PdDMh5t4LLvwpdCY8NInxuWdk/go2G+Xo8vA5cMV9cxiOxTaiDH/GxWuwi2fO6V4Gps+
1+7I2C/Y4doBUYDHrx/wLsPse7yeLc0d2/JGPBFwzgMhO2S2rm8UxJ9OIZqp8YoJU8cjtsrf2UZ3
C5gIyVi8+tqn0KykBjRB3QyO08l7KibIvyXHC+pYuDkP/oH0pGD9O2Dxw6ZAGd/jOt9JTZtNUt5J
Jm1VwKBopsW9cMP3F8xN33z7H57j37LplYnxERiM3DoGZhexrCi1QFulOufRAZSkZaB+xG65VAW4
rG/vokrZf4qvuMh2d6dfRDuWZC1Ac3yyvVKzIUzhe3MiBaXq54Yj/Fc0zhmEzwiY70xDMHWZWo41
i1y8sJIXu3qr3L9VTRO/wsj+p3NyErXEEch6HbCR4Q5mVzLhckmECRDxVfVGp+4j909kKL9E6/vB
+lkeLPYNXavMFEGK6toLYU0wslcdkh8o6AUKPyozD8398vVqozN9PoaYJm6OZrt2e6vNho8w+GID
S6C/FolpPSnV5M+hj8a0myQgIYpXExEGESt6YukJbMa+WDk24BCPf/pYj2VwQUf1o9iRDOwn0RA0
v7m7RW3uh+EB18kmJNNfZqJgIo7uIw2s0iQNGZsT/B1bG/nYPHotEUUxktlKipyRLbrC8AuKXcET
xKiXA894MKo0RWopTRDXdVknQagOZDmai91Z5QOtaI029jrQEfebrC0vTtJkOkAo/Ao4v0tk3eRR
HM8XfmYr37JSKkLsZh/Xp8VdhKCJfnlnWdjQyFYXCwGVPRSHuvdQauW/KFkdL1GsE8P01eEnYTkm
fUsjtepWaZLRfQ6euVSAsmolZPbLCu2hCITPFI2Fty6+WTtaPWVBRRkG2GsFKJAOF7uM+iYPsI0Q
XTYOn4geI6qSZZz8U3GhyIzb3xv4NNjUgQIVwkM77tgkh2WV9mK8aJiYXeUGV+zd76SZisK9TgMw
gwUY5dGbHHL1/pDPtLVBbd2ekVgy3+0EhW+/HVV9MDdQxfQGt8Sn0ZRqiB/POoHQWbwlS0RkKMXH
nC7iYz86TFYp9vONiDiidAQSkdfCD50mUPXptZN/k8iJaOluWj/1LLuggmbYxzMSh19gQpd0wtez
1aKDhAW7DxHEd6AvQrTNzIi99i4kak4OINR8UmO9r13CqtFVouR2W2QvNFsMTzWt2XAqec3w9q0I
gXsLtWvNFKydCciLzipVsw88Vrc20x/+4DS3aZVVFuvG245e0piqA2rJ8eHu8dLMcMrYkAaRu970
IIKLn9paAyWIbzMGoOJCOxMxYYE83FTPHVWk4LI6HOOtIizbJNb/tindhVuyo9rQK6l0KPFXA257
GHcPVbTFcOt4Rgs4laD79WkMgrVpvC3s56fmtrnCnaB7xGtKlY8+YxERbToIeXE120BK66l4AD+b
FAYXmPsFN/XA7PbiFuA6iRWzpq54tPGBioX4kkhwE0fwRTXS5iw+LUn/7eEadg0yLKv1nFIP9QLO
SyciEhMsivdMN4GzDXWqxr00kW+Qbkl6GJssnvR2IAmgO0W8kgYwGwTiEg7JGgK15na9aBM/TPd8
fZmKg3IwQE00PblrGKvP18TDeWoYDFOyz2gmR/huatPsjzhKLJIhJtAdAGAS9QbR+kXKbvZipO5x
1LVEAwP548aWy2o55UN3ybCG7BAHTKklLWxw27DJI4D/VV8L3dSIFAXUyvQtqteIW1xbAXtRfNvQ
IqXPa2ITJpfmQYvZPD751FcfRU/rfrOmMTRenwxo+/7Bd5PCfc5bvRL+63IeLZj83pFTDZuQY8RY
7Wt6OXaoA+HvcFO31srx5Ce8U8m67MajuSvD6Vr4c7Epe134isaWHFnJYltDE0ZmDNyaGo6P9Hxl
Yf8E+ZLI14f/HORat/iMo2LvA2dB9fbkJMPEcoCeufy+U6b3K23yQQbYEh5piTRCMb/A+hEehkuI
JzyVBuPBA9oOCGVze6aZE+kwPwDiYMvvhfOUoI24n2WICCqvXPEOR1XsNeU1S6KRjR4O74OnsBy7
23MAPMlesGwxQfnm7OWQ3pvSkETGzYpwSEBeek7TiqAu9ti/QNb0V6T/GbbIFI3HJL2xjwg5Uptj
rk2j6iVfWwT0OABIbInFFkRMKCZbakFLlRZY5yOoUpP1xpoLir6BRtXD9Pf9xwAPXzx5b5R9qPCD
s0usMaiD7LDbFo1V6Gng3SVEJ8c6OotioFD0lJG5G6wi+J6sCP1DjTDl/lvpiMw3taTQ9VwmQ+Ta
3M9y54TuCU8kxwPtA8Z5zejK+bKKb77VdOTF2+0AnKEnba8xKQwVBnB8M6TNGuTMhUynxmvlOQCv
erSpI8LQhNXhl5QDtfDv6yrWo2JUGKBolNPE6Z6ZmW57KPcrplrPXS2RwnRC/efcniKhL/v5F9ya
o5ulfxf4nbflh6XWvxsRXs5nLPEeub8vqsUNNr8JJrgMxldCKoOVc4d2i+a1RJM1B0vYk2KRtCp+
eG1MPcIuHkJe3sH1VRw5b12mfimGn6usEPT5V8Tm1W6QCUcxUu/XZoroNA+aiPEyCKcRXs4Zd+WE
uI7we4uVhPLS/zBVgfeHsy9wmzk+3YAjHkzd0BdHWvFifk7wTxhNmIFMSOWS5ZqQOAU2KSiwdorK
RjhFQwAv9xmSStVvM5iMR/plGASdOQPGWy0Bbjfj1T8elS9TmS+VEdkU9gHPnCLyPArpSoJ+h3G3
SK/XADEQQyS2zMGHhN1tDtj2cEfPI6eATYlDdbFScjMjyv3LKhNmTy3eK24fnrsUO1K9xY7o5VMK
EybYkLajsBqqmi/xAo24SrSi8Vobd4HsGgQku/5KQnar9wk5t0t0kjoKzjGXyH9AimC/p4jfKD+g
16ZY7kGlecyaXyKuIL/gotuz47YO1r34yy8/C/N+lFzhcZFPJqPd31AfWeJuVoCVvBuMOSr1lSeR
S69J4403a3VVKBuL2jaVJWs1hwaQ8JzLG7WeEoURsKIyAwzDmv92kgEKBl/MkXRzto5WkzGGbqrX
Mom94RcRefF/nBDzcMajUVxC/fFpNtHHxDwanO6zCFQkeDmghd+TnjWflDTHOiZtpnIoKuBRbwaT
prga/GiUL6ZdfLVaRR3qXqrEYQ97CHd484k1m94UQT1CkcwBpyIq661lanwLkr8q3V4xImtRPnlK
kTeWJrTKeeLGSs5XhbFTiXlRp4ZU6+xgZxBTdOstbBMyDp1OnXFaMuvTSsSR20VYyZKXhw8VkVTo
HAUGf6DF5ddl044wgX2SUoxOdQ/XIPUpmZuFWyVvq221F4kMWcalsgQQPvz92l2oj7PfafcpacRB
UXCJhFJRoUROZRvRA+cOLu4DV1sj4ukqVkNMkeNDxgL3I7yQQRykJabTyLtwClhCL3vff+8u0zf5
uHkXH0J/yIVjDPf6yVZvJwvlmvsjPpG9U1F/ZVNzOxGNYFyOIrTx642c63yFr7/2nipNNdftc/fD
VUJX+z0pk++l3NijIaicIuMvcX1k56NY/9EfC6RuWaGV/mMfc6TAMGhxyF3AVXLq4VVqTGYDQkoh
9rFivpVOeqzXNTsc3rnrzwCtAGkFAVm+/T5HgTPTXdEiVnvbUH5TNIqmXIz056/OxaSdixYFTpi4
rET6GrzMqvk00lnTQZaBfEfQmiJOwRZzm3qwzwf83hVFshNJNSyWu8SV3rhpB5kxP1E+5bLlqXRZ
S4higFzTODk1pVArwQme+OhFDPNfnhNUM1eEQs5h36wZtNFOwhrCaCBKDVXPZWQ3apkGh2k66l5u
lWm9L+S9p+TZOqxR1Y4ccWbS4bZMS7UybOkLLsCacubL2bAu0b5niLed26mzKi6SZRtOiRhLhoVm
X8bpczn4pvDC9r5DRcUhoZmC6x15DfIxZ6WNvKI0u6rYvj2PeTsBjgbQlyj6iD3Oz7nXht1C9dVa
vZ2id7GMjUzIFGzzPMBy0O15uobKHaAXfrI588y+a192QacYQ9cTsY9MYQwhf/qGEEmmz1L/R2i0
uU9jIltUrouv1HaQ61jKUs30I3CswVH0pVU+p0M5HHyPUAR4bzQ2fbifuFeVs4YP1gHAm1QVw+Cw
w/+GWd99O3kM7Eq4+MAC0REJFgYbb/EUEq8pwT8sJ/RiNoMTlUpucWFj7XLwJ+osCJOcZ2ktnLVD
xtssBjo8famxpvA5ohcVh1wEGsHEdNAdVhBbb6JBL+kQOYlitWPh0hhMrgkWJUzwf+UB2wOsbPZq
IPxqswnM4Fo+8bPuBLoAVWdXlfwUOQToV8uW2cwivLh97zYqSzjBlqALg9E+Z3Taej0+beV/S3h2
PqwKZ3ZPVUeRUa9b5tTRDDD7CFnwrD0H0YUGjgej92QDv3f21kM1NobNMh57bqN+vhqOXoCSVGIV
jKay3p/4fvTI3X+mJlzt7ES+Herf4o3mUHFknebEibecAgwU8/u8yOWeCjJ4MBH4o5tuxStUyxpr
By0Hn7+azH7IA8ChiCllXAyPGmyIJ2bajdp3dTJ/uyW1QB6U5zHLLOjLWHBfSZN/frm64+LzYu12
rirmcQgjQx30iyELHnX6NGCYmu1SX3CL00A8/B73gFDyrFGELzMoTBMzTmxSqLHG2ghse9O2xeTh
JemGd5F22YyVkdtHtPr/hc8VO4RxgxeO22TZluWq6D1XYsxXAPsOpXAZioS/ZTZag1Wo3hCZvbjr
8PovCUb98/kStnqOHehJrK5FVWFA/+7My2xlq6oqwlq6aCdXI00pmF8OUXuOb5FbBODpWL7cgTqI
d4pWQfmC3HUadAVWMah1PSUe3RjMqvVgxSc31a2i0Wjxfb7bEU8TWcNikE6FLelK208RCAWgFCTO
5r3jkxIKiez8h1sG8PcF0uDIXwixdZjT6HNd9sd4FVyviudxDu3W81diLuKcJ5oM6v3JMIbx/KjW
Lw/jtvCZR3v4mLVbz4VD7dy3PByaRPfFGxMYNI06KylD0sh88Iict7p1tacTLPiF4V9m8EHPynVN
cCP7u88HyozInk8KN8yhkVT2fzUiKyOhcIhzFunnZRf+IOB8m26NMujOV4JUAu9KkBlirPezZhti
dCE8d3zt+vhXRRpEQQwATLi3Lh9O6Sq8rQDQwoGiwKT1Yfs1+KS63uQWqOFWYLO9f0Rjt6nQl1HR
Uv5/qJZp2HSzacCLp+6BCt2dX/tTtFT81jRL6IraFt6SuO2xDma91sSbtrsGwUxKOp2XsSHUaVWN
FZtw5u7pxS8ret1WGAjof/gvmlm3/Qf+BxnMRB3M3S0P4KIzfr5rmfDEzEQdlB3rqGj4PPEBi6Cz
VW/IMFXWf5+jmxVOnbyrl73eEY2e9jpw2xyU6K9i5DlMX9J0AJYr0rRiPxyRl/fidF0EtQDmCanq
CoCIb5KX+UA2s5WmZVyYiW5/cVWTuktU73OkeF2KUWsOI828DxxgqGix8LOKtOMuSi7u+6IsYAPf
vhn2va1xTym4QRlNGjvAhrfp2l/DVuEinHJ7zcQYEwhlKMkLWdbMwGPBlJcXvrR05wKcOgZR30wE
8KdKH9sd4U3wzd2QXUjGlNTXh19vSKfr8YhAL7A2LKRZOUkQaXRBQVDj0X59IdrghFZl0b7Siese
M6YYqXmE5s/kUaMLNtIQSLHacxb5EqjE/euR443J+hr2RoC8wq9R2ZT0qayE3OPzb+M40X8ZEBkM
1pkBD5MpFCAKaAleIaHFBw8ysBZrSavcINKKDeHW5B3mXx3wZBhy4mZXiTZ5Bogc6zwpAMZLtLWL
9z4ETMINIbJ2yieKsHLnEeDQrmVXdLuCvkVcPDQr8w3n1Y8l/94MBZ0GOJW/A6TSirrZ1GYCu1sj
3Xws0ZtqMakULmcm4+Nhrx9K1jh1yNuPj/P/yAr2U3KyHmcO3BjYAibo4qwcdJvrRqHNkcsjWRk0
pXhMJZ49k62HnSgOH3axUGsnpK3/pf1dRHdpaS4DgS97b17ZbwgF+dTJ1/pjoq7urXDTppVB+yZ0
ke9tS+UXCLMFKbiZomY1YdupMWOeOVK5xSSVxt4kCZZYNUKiU+zityuqQzFKMtWfqbEGQ8HR5rpA
4K3pncjJHJVf8YSDihQr8SGadigIN2PxN4QYPzjy1QKFbc/m9MsdYhIZz/JhoG3pduxYQ3I+Q8Kn
K+FuOcFWLIV7gsxfNYfdQWiqquUK+mkkqzJ9Vkck86tiVCi2n+P3Q9csvbDYUR1rwcj30tgOOIe9
jFLk4nDIwVwDnp+8OcRSIOee/AgG9KVFeREN5Ajp/IIDXhlBu8xO08OHC/ZePjlHpJwHLtQhoYN+
uZrh5Nija1QzdQOnVhaTEEYil6xvk8UfrmGhI41DQIgMihC1fSbc6TXv/jgG7/pc26frdstkCTfq
9DCcbg75lZpEtssT1/CCFLy3o3VcRuVAxHZS37FIzLjVHF7gSUIlyPPwcHei7kNeOpnA6sX4vC+s
yRvCCPuOUnAfxePV8xEOP32ocQww2aQ32NUEpkzrZYrw8G2sFUugMOF0a8ZvZ5I/Z6MHmuTeJTuO
xfe4C/lFbc+3tfNDPS+SJDWwUcxNjVbWdhu2OOxvU0/6lUWBNXVwRrBSyEqGQLCCbOl4PAfFBBI4
n/3MwjHG5b9Xz8YmcDp3OqkmL3Z0tmZKEHU6XRjTXVCsRPD8196/gAhmKPOHWOrdq6hHD6ssMAM9
F1+ahoNrppooOc/3zpM9WprS41ifXKTJvaPGMuTx5r9ereqcQgtUtivGQ01fNLBPRIXRjAX2Aer4
5E/fr0TXS+DEE226Jg0sU3t0vsSNw69NJAIoj6bG4xU0axovEurLa+J3UHTUX0zaxFXFd2hNahTg
Yuy9Ugpi44ZCqUWxpGLPjI7TMudvnAUa01SGkusuJRAOQg1nUwJTQnMzJ2yQxuOFiFMA04TsEgwL
fWhavVRUVnWKVGOezVAnk1s9K03G7jmNyWYt5SZY54X+9SVjZEs/NPmUAHTP94LDRPsEmnsGWIou
S3jwMozWJWcoASt0xDx1H61BccP2zBLRl+AX/8yqVQ985jaDR1E37C/RueKSq2OWtYpp4u+nhHb7
nUjM0WIArpEcEtEy9x9TOO45IqhkzpxLnyNB3wzIVQXDcSMnF8ClRPiu5Xqoc7DwZ2XflgFQMLEd
nwL6gO2nYxSlyBWFfdIQfiwirq6w2YWhT29uGWqsJGsjCpSvEm9eYV/xvvEMJAFx4iUYGAGOPT3b
KpdkXG9cZsvFPhyUFKXjKbZ+boZfKkz6GtyJ209fseBQIOXC2jrGR0+az9k8J40gH5++X7Neantu
SZgm+mCSrhIQ0J+y+10kZHcxC1gWcdiHXOtnHgDqSmz4sMwNLP5PsBUu/JvG8tbClvxQejpzLGhw
/kfNsNX2xmFZZ4r5GnzsakkMOSrSqASOqBfDcyQr5hNDXA0DZ1vNMAldyBgpnAYwWdu+qmuPCpHf
LzG9NLDPaN42Ubcc9GexMURrqVcwWo/kUSyYf89ImTLIFtknd/pYsaR57Gif+unImSAgbc5HbzLe
forThQVO05LhvK41jTG6t/Q9vhE0LM3ipaWYlFitSGgZF7Ef1Xo90oDGAtp2aDlc1UnkvdnEPIkE
cDP7k1Uy/ZghmXe1JzkwA2YaA+WQu1dN2cwWc/j/xRXZnGb+vTEca9utaJc/sfmiMdGRUtv8amDx
tRYaVvBkrS5wJ5fHRY1F1WBABMdXbo1mMT8JAWiGYYkqpgcVGmo8zpm1aqpqB6Mt7e+WE0OjDz27
BY+eXIWerthiDUwQMLYUisMvxL15joQ0nTPKyLPScagmFevHdozoZs/8Vx2zzCRf+ty7xkpCUG/l
522dhzk0E8HNHZq3c9O2TL4TPMKmoitkZ81S5oFafjsq5gwCZTc4tKDRYDhpmNuGv5qlEe2Ezn+d
pkwQ9xOPnOfpHpPvOhTsHmhqvv6+8yryKAPPYUHtSUboYv/qU0T7iKvdzf3GVDX4Xphq10hvsECg
/Trt4D9XNO2Q9gY0krvm2dtIuYwdL0HmXHg+vBbOvkR5yEx1mXHUZGDImz/+mgTM0raRzuJ6k4hU
IIiHw678WmXyUIBfsE9VkuBLOOFa9ZZVQbiKgo56fMJ4xAXYHqNcZuvdTXVuLi39V6eEyjrKUB3S
gXvXRpuXtu2xl6IW0flJWkEEjVorb76yZBX7QmIuZwX9W/oIKYs0WYvP8Qd9RtIJLSCyKgbfvM2b
bSBcRknDSvR5FM/Afo8N4CbZ2PE/xUzbBkwbGCmDdq0Ch9z7b4/sdMf2eSADiuMFFZoybr/ISVH3
WDZTeMELh/Li1ODKPYR1CkpFjvq9QhiUzsjZD/3UTz7aS/dgX77jtGq260jy0LHVOz90YI/VPfD9
Yl8qeV4VHUNl3ewL92A+r756wa2BuVOcy0eSSnQ0MJeafNgHZjl+PoNhgilwLp3OGAJ306wElOGv
gQ5OUyPXA8OmyY7XAxu/xXlQaPptB8K3DiL4EN12IEResRVNeGYQP0vlB78H9mtgrwXGKL1E2P+7
rg0sgSQIDb01ewkdviSn56XxpX48Qjxn2xEgW4aSFwnGKvm0LeOb/wSe22LVipz2MQjTHbhPX/A3
kTcBsKwx3IfetKpDxci5f6UEoDBmGVTHWdXcCHUfY1kfK3GMR/gmqcMFhVCtO3Dv9YGB0xKsaMsm
LkP5M+P4G7xJNyme8Ajn2yiQnbCA+OqVPOECrws7hYOn45ymQxSENXVOapp2/wlDOPbMCjgQftR3
iXhA5+wVPgJnef5X9EJv5y8Ocvpom0/s+vkV2exDhmwUFoleRrKa7HfgGLy848MFpojMVgPDK1sK
gBzaKLNRwnL1vVpEeAtJNZ0An4LvQIT0QkBpVumPKYhLL1fRgeV3oMqJXfLUT3g/+/+wQq2d9xsk
PWlQXx2oJ85CtpJElX6Aj4+3T8HLF3ZZat1Mctm9w4Y+qzFXpvMx0GwcfzWOVrA7T9+U7LWLNAR6
q8XErMqCJQ/kJNbjFlnP00IUIDGcHRB/9QySz6dh8lQthK/gJ9yNh1kmSZ/agsWGa6HlxTnlARlO
bPb6MCerKnRxuA6TM8zS3mfPw9DiDKAULOM/fjuPkSzKhh5ERgkRP6YzVaRvQYrcJJ+9r6SdZEL2
YkdKQsbDRv09y3lMrK0een7ZyjAxgU2O/2/Y5bnpgN/xKjXB2CR0JincMg/3ByIUAvGTnSo09+UF
puURyw0oFQrby5yi5LlXzVMJCXzTPpbas5Yi9rXwPYBZhg1ctVIvJItTSXhrMq4jfIubZV1gb1SC
Wl4IGhqDr5ktrznyWhz6pB5Nhp3aNW2oIpC9RJ0E5lrNim1EJX07gvKrvKNQMXrfFpJYowNGm8Ik
KI/ZesiX1KDU1kY5LV9CqYvXPFsFqAt52IX7OmSbCwblS5fA7QOBd2J8LqA0jxMShpdRKvVCsTE6
Uz1SwRe8GnklIeAF2ngzsHFM5/N24QT4wWpaA2xeBKdXDo3ABhplWOo7lzFeiVQZjCaI9KOClatl
o9G9ZafCnjSOVUDwis1wuOgv3VCGlUWi6SNlQXvNZc/heJrh/XRdwNrtiE3SegIMSkN6Szm2Qht+
HvFQDHmFcCdMhgj3F3VoYqnxBxhi6mTIw+srS1ur/v/WrqcWfI/22l/gsDxHHKs9tPvy09iljz5a
/AbrbrUdD8bhGvzgD3gUYyMyKsaVGL1OlTuZLOkL1jdLOPuUEpEnnUwGzaxt7U18XspMvTMeXvAw
Kz6nyC4Y1Faq6XrAPuF4YWSkg/eKiwE/NXMMZhhNrOpYqfB1niuj1Hkkt+NSTRgVqJacGflsbVvf
sepZhEeVxzUDbHHCKRII0bSo+gk4p1RcZlhR08DArcfUdlaCd78jN25Lvxb9HSYG830DdkLwPWOS
fcQ/6OAYL+1WQM/HPO698oU5rJBMCpLhVKeC+5va852tSSH9egzFkMWkzvWVSO7PDT4YzlkbZEeA
jyLkZ37jg0aDICJsA8Z7TE54m+pmxzNxh0LPzPbd6NGvjg0YT/OW8ZbYdFdNAXKzqi4qyvYWQ/MG
vBLB3GYaEWLJcgsY6obxalKUKQdYtPqlu+Pg1knc//Ihi4egZGeqb/nJRwdiken0sm7t0yTs2lei
AdWRvjhD2Sy9xf0wdYdvBKej+vJS88jMxwiaV5JWsFL/ZQPl1vQf8JIwFPX4otbnJZ+xtkn6UKXR
wJcHa4uBkOmGp1Bl+q4+S+YADd8Ay5eObJyAtT+afg4xeRXfWeKmlTsCVkEGQyi7u3ULH1OzYsw7
HP9xF8oaxWFPffpoYJWhhUXiPc0YanxeXGC+o2Cny6yG8AFXxOngaA3Oz1TZ+ssbrsDFNuQn876t
9l7l9j7DvucNsHMb4YNI+KG05wajLmt6iex0DhAdXbH9wy1/XBifRzLBzUpIlkuSSxrD4PBiWrvF
DviZJ2MSP4JKHP22fSB4YpKUDUkilVW5I1iNvE7PmXGbAehQhhBOF8UKDjdeDF2FJgAYfO+78yK7
B8JL1ujdXL+ZtOJLs35rmyIWMzOEaRECilcKXeiXi54Ig/fDOo4QZaNb/R9CJ80v0My6YpeQnag0
Ka2kSdSvvua6ScqAX5RuybUesOD+qK5v4jdrWKoOcfN2oru5MLMkJ79eY7MFMgdD/gPj5MdCMPmd
EGYMOa61zxMUNXkw+H5yseEE+4XE9nmrzgWlcOekYrVjQSN1TevKCoUTtPPvVNJJOp01ND6KXS5H
uOSxiP1K/64/bvF0V/zkqjBF9O0hlHRevu3uHNVyKDD30joihqklZ9TXxxsHr4IHbbXFSu7bCaR2
sQBiQuoOK0eMjzvT/5q2Si1yTWhUybvfKakE2ybLqoKu2BfLvhpOOGR/wCdyiiTUwb8xBdvHfEVX
ummAKjzfEk7VXjZIebkhjG+MK5sAlERkR+woO0Uabps2qanY2tyalZ7zMum0Wmd74XSuOsI7qne5
HDviDxN/0sRmhULrxEEJHw3e4/MGzINUE2ycmZvEP/aZ8iSQEd94drtSaJ6Vak7g0wBFfAl7ovWN
QCoD1Y3sE0Os0S0mkVPGU4Pp/UMDt4+1uH4cOA2l6qVoEJdqr9JXTv6/59gLRPoHFBgmAtIQJcNU
P4Gu9PSxVe1lOlGZeu802aN8Deff8KFl+0d3yaokRffzyiEsWcEYpGuH85aGxaBlqPoU2P9Ymf2U
q4cbabAGn42Mi2BpieE7uPfJ8zt6lFqBXPi/r6xu2O/7G9wqdYr04hp1iAxIEXlnFY+nNd0MZIDj
1+mV9Vbk50w0p/c/Qy6V6qPfQK38Q+QXBwkPJKxgwrkKZH1XLPLkw8q3p4ipVn4swgQLIaRUJwAz
wyAGdZqq+f/+QIK6wlREo9h2rf6wxThTXhukSLovhkN2a5dDFkj9bZPWES27xTLcb1NRPWbr/qRR
leD7p3EfAfI+VRAbTjGgnMx38V0EKbW7MF6IsgKCMJ0QHE3ijlsxJzxfHuvfoU5KcHJ1EVPCFS5K
miqCxd6L4GNbtZxKtDltGgYSDyNHM8U5zjoFQzEbE89dYn64A5La1iqIlhru29Iwip95/1goWlxm
KLY6eytrJD1ZOMPw+eKDJXeJRLpcqWirhI2V0tuRyiw/OROgp+j6M+1oPkR0Lc0VUeuSzt083TOP
arxCdsdNsy+nayNzIgazprBaOE7GNZqzj5A02FMGT7D15EY9guZshLpr4FCsXlOeIdtAbut4G1hD
1UaZ1WUD2VCvGGy5jCpJGQUSSMF6e5glhlydA794OTfhxy7mWMVfRDwgnImN5JyfFVmDPubvdd4t
Gaai9ADhs+HPG8SvSpf8bsHaSbqGP05WvIeSSWWF2BZhA5iWPkDpmS47UvE8lm7W39UvjtjBiS6S
5FvYFy04Y1rTh21pJRcSSLD934asCQSIy/BfHBQYzU9XAMspLz13F2T78PWQh8//1io11dhQ3g/F
zbJflS5ghBQDDPiUl2gauQJZxRIURGKatcj7uysWLLBzfEXDTGhWEYALYhqz/1SNrYiS5I6B2Lt4
GTBBnric+MAhJo0HCHU8yMjk5EI24GQlKaAC3m+ljBfGsBDeuPUbv/1wmbrrQ5pc+Y2wXrg3G9B/
z+bPtwbk2uoXleUnzgbUb7cGUxBIK4U68cpwykgMoDcPeCotyhu+CVxcgi2tXnmf6rUqSEGtp83d
qr6O5zhffc/8z7ULExZ8aIKQhgvpjWa5964A3vGQAm4ku0RWsTdXO1uJq+PbXVqoWafZ2if7GYDS
cuC8BdAhO9hXOnHLMPTveUsNu3z30TLxbav/1uB6HwT5IDD2a4Ei253XEu7hH7cBCTl5+owqGcak
RLDBWrWw4O1aLbSBzd6FF88JUunyn+OodmJfZpGwpMll5LXLuEUs9xe/OdRbDyQKNQp16Ls3x2i+
EyEqNuVvUm6WpPBXEqkTTbeROanr43AVR/MWTMH26oK9vK38h+Y2HvCA7y7jHS9c3xOh4KPvJxlA
6ks7iPKQxfEtoM3Z3URydFCv14SJqZKRzLfKMBE7xsOQcOMGKJFpfoMKmnhXBCJrRE+q0EIsVEDJ
BOhc+3+8dcCn1IXR/urfzwiSdHFIhBHYgBwx8xHKzVFpUFAjlMulpyj3yf0LcP9K7qxYybKC26hN
8+9ob/X7FG4G99rKelH7Di9VWdxppR7D8mfrssIwW37pkA7FFcQCI2hzMy6x+dgkVRm8neujliad
b9iH1r9tgbApFKTKyXO4jgJ5O2BWYxcq5LcJZzMNQFdhBqUzZN80lcpRKRb1rNRM2EVxHciEM780
nhitk08ch3R5o65RM4y8RZUIB4sCzZkFcHuRNTmHeLnUn2U5AtAsbcNdaZeJNK0n/eCuI3we2RP6
OPk1+ZBQxLInPDuIlg9AS9tl/4uxIdKc9HVnPgEWkYQXRdLJOaXgPmVgHbY2kAGI6xthV/N647MZ
gp9OF7eGIlogF473f078O0U86EFGAn3/fVCALHujOWInZmy9X8dQpVUFI6abDKlTNjqLR7einxdB
K039GuXwAi44s5lyVAze+sVFgljWzkSIneWj0zxL9tP+7uRhiDj5MVBhPNCZT7UgTOFtNEd92H5W
HH+NBLmEPQZQtdK4E3fRJS+x3G5pOQKdBzIx0FPW5C2C85oWuwCk6pN6l0VJFSutdm9jGEJz+waz
x+Eknbm4pWABffCzEGbe4elQ7VVwPQCTIM5OkQ2pDif7uPOxwZmTyC0UXFjo8Olp1nSlzM29uPZY
sfmOjow5Y2B0MEh8kx4iRJmNzr+UShOljjIjDiJMnMQ3i1DwI3VgXrwQ3dbNqgMOzBySjHQ7xwVD
RiOeznUZdYbBs5+yiQQddnjFesbDxow4ttwKSXc8m9zUQl5SKQv+802WWl4l3e/fsR31oHNTTuWh
+LDzmBs538Cj2cgCR7s0AJxz8OJDMv4FL74T8rYDUIEIGkV73K1ub1HbHJZoLN+K0BMR+3uTkuLQ
TwsXjupVTU7HH+ZpHl7mopw1c2tr1wSv6hIWuGmiHQpDuRO9W2ZAgJzZAvZKpBm+DkapfgRD0BeR
kzgaXPh2SeWRxbgMWECuqq/oVda3gTGTbjyt1m7nBxDVvJa32Xz0GPA53oklOZJzK4yn3FslGLn2
81Sy0upnNtukKAxEMjpeC6FJSrqAS/HDipgS4CFNlMVAUkkh6fWgLdPN3vcctmhLdI0IDkjit9Jb
nEfBpsLO11QrLGaqw+AdA8y+sF+SL9gjOy9csiUjNUmxByd+1Ni1nr8BxCKXUeD22yJ2xvNealW2
hP9TixxULWYIPw6lUFeiH71gDkMww2W4oFyVkA7B3MUZX0YOpz0iI2nqHIhGgWpMzGlC/rWY3xin
y67d9WwjySI7qcmLvlszAqGOUYwn9IgeJbRJ+uFgTb25uwAAOWeuuwt/SbY62JTLN43USMJq70lf
tIFNRlFjucQLVuhr6Su+2U2GZq9g0E7lPsY3wznPyPFFxwC2UzCDapY4vVMG2KKcJhp6AFGQ22zc
B30Taygnz3NRixmJi/2XjLsgZUrC5Of13NvUJ5U7MVSTQN9jbIPj1VD9ZuIuGwCyE9r9+WsyLsLV
vqazjxeT9h3R0XZfo9b6Ax3Vp7GXOeVlEFB/eviGFa1jqTXWsjSB48vyWR6LJ7fiTzaMj9vh7KL5
jRP+QCNR+GLgs0OkIpOXD//P8FdJk8xQOlXcaDqMVSw0BJAsyvMEVqEwsvi7PNLgl+UvMqjhA37F
97LJsGE2E9StBldagEtR5dAYiCgX5IiYQm59/w1ZhNa5evMDZYdc2TwzLltd+zcGoSqRHZW/X8Fj
Pz5nXp4ukV9q5WbuS2a5lrN9C/asuLJq5IJs+Asbi9BW+58ce+Q1TTvnNJyUqKJDBvaFouJ8vNtg
hz8mYpKst3fV7aziTZYq8HTbnV0IVW70T1xR9L5f5wmdkfRR4Xqtbl4JoYY0uIBGmmYBdVH2SpYK
h/Q9O8k0rPrKKj5wdD/3J5CJFxK/0whu2jGiHXdXzqCdJ7uUrnK0bVcVkl1FtgEgKkGzxDSCgn1p
m08kuWCls3Q6LSNpOsvMlJB3SYrBF2VaAZyEsXOrz2yyxMR0t8P+fYSYuCa10fW+Ogq4ptcIX5Mu
OUyHrhMPHGB8fHP2nz0nG86+Fq2niNUZvjHVmRK36Kex4y+NqWU/j6oG+XnZmy34SkyysdLeGDuI
ELK2wwjGs2N5VEvnHGGFw20qTSgQhIHR4QEgtLM8swQ2NU0riE57hLj/1FHDppTaPMV0FuaYhx7o
145QoaLd3AZRxYVzUrpNnPIvnQKQa783z30MEZEput6nY3ITBNE96OHbhVVmz7h8kDgvQNM1cdHf
hSn4dYWJ0qJlYvhDOk7Do+5Iqt0utKojaWnus6jDpj1mPwmlekPFlov0sLdbWKBrs1XhJ5lDF2l5
9pAEeD9CcqMFkpTyIdFcn3Aklv5b/ERXOpMgD+i721uGdRIYNg8sNxmwxzA70Z7PWYyz63Xni2Oe
GWyj1lVB0mvQ3q0hggS+r7MMkwQVaA/e/sV0jDgwN+SaADNOf8VYMkggyfrfLN6kNz6oyUpVC8ji
3uUQHJLYZuTjwGnDmd6N+YLZ6RIurHhIIE4y4+/WUs/5FX8DBUgfW7BSiasgLfyMqpGH7Y8Rgr4G
FLAY7wORC9lpMqzKbT5I9vY2MUxg5LKG9l5BA/eEXLoo+JljeIexRdj2f3yFQEeFlsUHlwPixWbR
C00EBd7feVOAHL4dEFtZlLsjapBRlSyfLfE8MyOBDzRKfsU9QTfgqyCXt10ulQRttY8NtAcohVMW
zAetDm5TNGIL7dxgovciJEN3zEd4nNiCFLU1J2HySfm2SAPdT5znm0BjVf7wylFvbkAhyxJslKGO
H05MdqwdAojxi1jMnyKVAlgw7RDmRah7/XWAU1UgSVJ4GohbTzfxp6sC3ZSVR0zSKF5NKtTpfElT
vAOG0WPoBgPESE3bfYygFYOetpgkBPuabYMYTQrcg/eFt+T7tDcHy0zAvTclnCBdxtV1zVujlbms
9LLBXTnyt1h6CudZWZBCknIk0jNUz1X+S3faL1ayoMte6CKbNKjvLy0nvKgkOxVFDdrOQjir9yc0
fQ+2T4Eo38znAp+uF5UMUExVDGCmrFYbV4WwyL4JAF/ckrNkNCCdy/11Iak/xYc9LHFVQ63Oy2XR
rLq67ZnPAXJxYFIrM8eACPlHSMdxp6XP0Ly5m4zynEHIqVasIYFAy8j9+1KlWrdb7+uX/M9sjd9g
GOouT9V50Iwa9A2Ny/YlABRW6GYFVWWH7DgU+4w7Y/DHhUHt4ZbXrHa303jLb38FtkaMNlqii/DM
EXyM078KiUyW3ItI+6O//u3YnF636r76kYbQS/BER2fKRkaZajhu21rI9k46YAYjdxhiqaaHEjzJ
Cg6pk4f7h1fthqLVXdorCL1s2Bgowy1gn9RJetQrrT1LCZXh9zkz3qQNGM7odMMmw5X3jXogwaS6
IDJjH8ulCbfQva7IKK0NF19R+LS/a2n5u8kF3AlBVO2/lsmRLHjfMi9QGydv3U8MTKZoXoyM9GYO
rPeEHWc49NUwlm7/6/0YiPyjllC8xfmV87mWn0KeSrIGBu05+9psuXAVMYdgX/cH02j07MFM/egZ
g7MCA8pD7l4JalxBC5Z3D9A7R48ZcZ0XgekENh4/PswGpDJl2MaRDTDUyeE5honNfp41YhS4idqO
o1pJqva+bVBCzpg8KnnOc0+MI+FjiKGxX1i9eSN1i7ID+sjDOokPdlFW9DDKyFwuV2cjIiU2dGCU
f26WkDXY1QhC6nRCJHQYcrsyX0vMRFBCRSVpv5XTbulux2bk21DibnZ4c/SGLNwYEi4yqntWcdGj
Lj6hoWcdnwGb9MiQ/8HlhSHs1iCGpQhTtmQ2n8+esI9/QLMlKBsoOKMG0om3J/eBVshO0KhwP8RO
hwO2YuPKiJHOXwG2Dy3CpxMWwqEy1XJ14mVkt82IVOuSgescB+O2LA2WMggbPwkmKMAWv2uLWM13
5CIQwCBtNJpJoS/fY9vWZHAlU5ySWKGEPYnqrlt+ULg4JnOXblW56AXRuLdfiSDLbXd19x6UquFq
L+WJK1pBFnX4yySz+2IJvE8jD1gfHyYHXNUIXzBnKFBx4ZtUEom23m+9fHAfS6Pbs7P/e24uPBFk
HcdNQzmtk7zm23CUICTn18+x1wdtOw1RWB0NtuKEGhveIdfV66xF2e56K3hVZb32nayiGX1A4rhV
oEgDcwZ3GxDSKUrAh046D2ZuAi+llKc9QtUBq+7NDIS+4K5BaQOdSCw6F7+KL8UGsq9eMwV7TvVF
TYX3TbH+HdIJfb1NNYvN1H6NH6HmEspovEP0oPa9abkLYM/v5zOF/GcmKneXY6+/wZeutOjCCx2V
iZy9AkCB5bXqHW2QbW2uorNTOunYsHJPFEw+BNBj4mx1M2bJbBDfDwSC0VtrirHQ8bhcJ3PNSCWy
WcMa5ee087U0+pRJrWiW5GQGX7JAM6BrdM7rMSP2idc2TLwvhmDe19E93lgw1V4+fGWft5nIy9J/
mQQiKk8HWqTQanP5vqkn4Oq0YNZV49XQTNatgnnujboubkxJLqLgj0r6GXF0+Cx6XqnqqWl4hHIi
91r5BAX238r/MnwsdleZdeidEuVEgTV5P0FNTkjr3WN+QWU6QaCZWTFNelijchRmqtDKM5mgGIj3
SbvhNYscGGHW17AhqFaXEBLpUlGwAgzYvPXfsvTCaJqL967J1OTxpDSlQVNUGJVlrZTDOzmPrFEr
h0cgBL73+gXrY6ThlzQROK9gve2ku51mTz/ufzIFsskme3NzTDEeauK0E0Is0jVu80mMHA5eOBsg
twK7tE/BuSbtLSnBoQ2WQzucC3fq6OyHl7WVPTBETKcwLXuinVKtOXJhy6TSBa6/w8XXaqdb6zsx
XPGxikZdjhGoXzhPEsntbBofxh46C3VQijGBbo77SOjbW9bWEhkgtzURrOY+HtKnD1w/QK4sfcQB
ZtWu1CyhIasXp7T+Am01GBhzfioVfTEeixU8q8xQONwfvKQhKBPBE89/XYxGfDwI5Cj30V9lFQGX
CVb1CvrsAGjsxtYa34VvJg61zuWFnter+S2zZpEpdIT1xgA2UjNJ5tC6FJya2S4CVTT6NAmVOa1V
fl2Yz3AXofgXFKQam0qbp0iezQJ3rTm4kY6WDgHlDjPcM+HkrLCsQROOx9a+sy5BQ/qfqugE+oBe
/3L8OyhM9JnLeDuWNkgt6MsGFAIvNXI87/wYCLMmygAdvCGYVIwZRPMNxVkKKlP8J74R9dRNQJmI
1XwNpdmMGbFJ+cf8ZiyJK6BssM8ky4Hu37GEWzIa5jqjNHLFSVDKHs+QX0x98ebnPncak5+jFSwf
ka/KrsVnwIz7DCh8XWKOhx3eOy5rhohx8XH/JtSO76KX6t3B7osjNe8XR9QG88XntG97OW5SMk15
Q5r0J7R8PlEth5/x5XSH5w+eB5mNsprV0mUQZp3WVTltkuc8ArN0e3ZUsQBccPmiCheudZHV3mvN
Svo+jljsbWxcwibmT0xSRDA6iddkTxr5tafPxL7YxHFaIipQ8Swz35dSrSz5p1Ctqd9ANVf3JzX7
RJiOejbc6wO14spl5arYHPtMNMvwS4EP2c83PJIALQKPCReUOUeeVUIawRF3Bt/G3zfRlSHsjmMe
sz80C2KTuJ207sxw/y5dbbeii+uxWd03VCinKQWLuMHuGBweUy1mdx2pKNNHNW+CUddnPKLKz3Uz
VTAytbJGNrv1XkpdK5eQQ8U1giT3kI+DZ5HYaNJst2FgJhhXbxF1Er/8IY2mTIwvK3uvnj+2eXUX
xs1zXUbqLypz9D1dFxC4U+sVidPgEADLH7/n1qB9NfX0/Sn48fGTBfyDlbe0WTRjCk9B6PqSlGNR
LYTtPzxYL1CuVnLCoqagK4Wze5zakbbG6CNPHtwAA0VyqHeqHbVxW0LzQr6iKGq+s3Il0NK5QZDo
ZK2r9onHGXpCkUBD5JrO58AMmvhd0eTr1WJvR05MqixeUlsilmuSwWjOCtsuQUhDbD/+8Y7cF92C
V5OzyGlmur7KdA0gQpmt3e3sbpUjg0XORh3Sffu5rr7mDb9l/MhGYKHguBkXeFqTB98C9MgvWgWJ
5gz4quoblMLjw/t/+4KNNrYMxLTEOtPri6H4dreBUZaMhE1X8cFTYYrug+JiOnTMYXgdyWTFZoSO
o3LrwX3GJTHYsg4uxqEHYrNw3iJiYpCb0MrGyxSeTjSEz4e+DJgH5cz7sy9c4peibPA2PkTw7JSo
Rylax5LP03D4AW9Wr1mzermVFKaGxhtslMiBmR66bGsrg5KHTuKITIogUCcNa8BkFEDF/SurQ/4o
U8+ObFRYTyURhDfkaSN/vq8KcfagNOmrb1VEQ2Y7U83+lp9bgNdPEV9eFJgKsueukxJNxYSgRvJ9
ZQFGZrAj6R/Rlw6fcCm3r0ZnFZFgZVuBbkAkG7Vp1niKKk+RVkqZiGHtb+RDcCJDI7G4/JiVPXTY
PBvldfiw+eqozY+DwiQ19ARweM2SfA7qxVad69XYD4bOTXA9em5gSInrmy0uVzIPATqoP5tYKaHc
W6n7LD1ZDSsBASEyZZllx6cH8tXzn4HPUG2JttwZCiraj8GD1wVmpBa9g+9txtIaU0MqezSIk6ew
q3FDbK5z/OumC+cTiaifoyufXwkXxnzxuwB1Pnc7ZISeJ1y3JLk+Ok9eD5zberYk6QU1Q7+kzS9D
YBDpgNVvjIPD5OZZJNfTiKHoZCZ2fmJC1iWpuuCxO6H7zP3TujLRmUwOQW4+UKQNEZLFyz6x6bor
2Sxfi4p7jME6o7LglcPuHBfcAoj4wNcz4F8DGRu4+AQxHGyB0WLEoyHhvI/ksD4NqMS/OGYYKLU+
mm7sOFIecsCOsGVfI43Azf8fIVkJ3jd6s/cioEMIbh7ATnih+IjVELqFVFx1m+nGHWFBE4KeygtA
gGZefQzOMLry9lqMPEUyfcNX/iTezcAIPJu6dnFHVFSknOP+vFPSEK4sZm/EIUCwalKt14WMpc9v
TxnpzokD1VZtttg7xZYgtB7FmNKKKaWG4EOaW+0QQbzllJXfVHYRPpQTRC3Q704TvzZhun5ZkAoK
keuFEqkb72WgmsxbK5Nour+R2N6oF+MwDcpxXH4FNuroJ77+15f4IfRRb48sdSltaIb++FL+ObHL
6FUJHFCHmzrRe2D8KX6JfmwtpdePe3boMhSt3NecG4XIugp5tZI31dDRXdbxC+KNJhwV7D9hs5yV
Pw9V8B852KZUG0yEQPxihQmRYmMV9iFw0utV2rOaDx6Euckneawbv3+s4r6hOnJ8UtlxE6oDk7la
jgCLY0OYd+1YbKDNwXSS0Rk7BZ0y+beSOHpDH45vjZ/TNT5aG2Qy6ZNQuzw9kVPtLGFmngJ4whxa
aFCymUcjYphUED3KiCd+7IJ/MPnR/z906bA2dDuuQdkl8SY52Ni6NmU7HCtmT/xKLJWVRL0SnDTF
3Y0ZxkL4G/bQzRVgHhW+2aaP0SRD0nnlh3/G0J2wQ9/drurG0n5QZkoZLDSfduNSPf8ZHgiq9UsQ
7tioK6a0KH+o0QaKEzK7Hp6fjODB5O/sgXwYYekh876QL2vANdVRR3HhHCqcZuiUN2NugI21Q42C
IVqJW6uaPeaU2gcPKx5J+3xn7YSUk1SJq81v0hTxo3vDl1HSwiwtiWQj0et1Cu8nOt1gQwD3x9nc
bfkmWpnGHDLzHIMtf2GDfbWvWcFVKq/8CjJGdmMDzOa7BMt3oX/mpah5+nRxiBKt4n56k9ty1XGJ
52+Uxy1TN19nZ/S2KOR2rnwRFxT4LtAfdTCHvzkhfzhzG8OCBze28tT18MY4lUTpaPQspPZVNML6
FfYW/+oST9MbUZfBI8TFwBnGUuYrELLs+zH10bx2W2+rrRtK/PcqzrQrajzxNuEq6wZdeoUejsmz
Y+iJfC1NImT/hnHukby4aK8mPrLQFAZguiz83hGwWH7ftkaSPMKRJqppN82tpIV9ApsQzCNOgar8
JRnfIOiLra74YdE1OjdPf6j3Ogki0Ybbwbs+pqSsBgW/nuG0Es/Iui5MpcnrOiRj3YBykDRxVGA8
WwhZnZOWK7Z5NoZ84idfTxaDKvKTCbRCzTpyzMkQUK1g9vvB5V+6/yjT4Nw7bMJiOGx30bToBEO6
FBjMKTzlF6QFSZNt6fF+qyIeuj62RXOPiLZJmiYpPgfVL2V4G6CNYvw6OA39ffV8yQtgitl48+yk
p7Yz/UO+K+sfQbxcxc2/7ok8dVEt3XZKaLmmP6/BR5tSjgPT27ISbDDsT7CEOk/D0dxLjyiEnu+5
8yDmUbNf7R40QV39eD2zQzRGp909w3tqEzpq0gsqaMhJGMRPYE7ANOHhYDPJJu6gUt9M7rqdtrV4
a1wBpyQ85l7V/ULrDxOQyFR5HCnJ/NNDSB1M2LzNasJ46CW62o7PAIeH/vMidOBb49kzMmv1OBnW
t04PfcYcnDwpynpR6F59yL1UPmZy9m/y3DChvQI4ojDpfjxCTJh49VAUXpvEg3zwPGokzVBlokwj
JwxAmaI+8W5+fqkiBODRu8jUItV1YWgYnwBLW8MbWXkLqY1NA3QynXXjjT59cyfCxjKAZK4mH2me
LbuFNdvM8LWpEWtv/Euen3rq2imsiWxcGNBoDBXcsKPenmzVoUfQDGKcTalgmI3IUZZjgBHmYbUb
xZfvEUZfIs3bKsyG0/U6V8JaBVBfSm9fbGz0sXgER/PT26PPSg5Ev57gJw7gZwie2EpWPoKI75EN
8mWM8+pNImVE6jd7fvSINBgigoZktBwVzwguUITgmH87ExYkDmN33dls7u9D3K0zMrqqFQmn8wbY
NFYKKMKthimFeeY+2i2i6V0ttQt7ifK+8YRlfATTLnkjJHwQc5a3icPzqvRmMwnnhqEgd9dMJCha
/Tu1Gs9ZxlKDDhX78Zn6Iul3ITarRUPinLiPaus0wtlGsZ51KRUVq+BkccD/3uuyZT386He4wYuP
3aTzyyHzic5E2hQFdO2ZpXnl5pEVis2p+v7/SExoecpNf8zTlnKOv33jFDocZMDVPb1nT0shBAz0
Qf50QxgZlEryYMSEplhyCVncmrwiZ3vCexGDcYMRXnedHvuFzTsggzJ+PcrmShCjb8yrm4be37SW
XDq9DbGyupfWKQ9SwM4uLZQ4056bN9Vg5zdOYl8cMbc6HGEt7L3pdS9FAVflUYCRKNPyo7CmpFd/
Mjx9hS5Z/XeqY0IvpNpv8IOYPa27BHkkxL1zX4iWZlYZwzNMFyzKjNTOi/QbDo5giEH3OEnoH74s
wZYnW54E07uS5ItdjJcwOY3cUwFm+wHaKmCJyELTqloX2/LgAb2cWwZ1DDnoij4O23IO7Fqp9qta
y7Bbl2vG8XRiWbzntvX8gwMME88O53Qtg2naiQsrLOMP95qUEKjZsyS1izcUKDAyxokqossuR7/L
DopjAK9IzOSYG69h6D3a2ewaZnz1bSpqWlhxLA7MeYsKc1MqpqIsEN19el5nM3BsC7oD6axz2xX0
jDEh8GP2R4eBZPwR6Cs/oPfbP2IIQu11XWPPQy1yQSvBcfXUaCTVMQFjYvbY1749VvRk5mkteVAH
E5c/rH76vonlr8rMWR9KSQVuvOH60wmLOuq+IqbMfPlYiI4a3N+J+AlSspH9FFzFyM36tw+UBIAz
cNlS9F3d3ucwDT6WiqBb1lW40amFcMUvBfYFJUfSWGozeXnUUOoOuNY+vDv2/SZoXTG24X2ZZPZ/
uMa4semXB3DV0eC+Zj/M+lGSK55ZrpKZhQgfFwr6chsYnQU2IgmMp3GoxMdKhinSA8Dj0ElJ3WsA
zT1n9t12mhWPmG8dAHk7WquN6pY7xgp9yQQdhYm43YPOljwnepINacxyDfnp8PjKLdnE3p8JcI3L
yTBWRXtOz2ceOJT/8Av0PHjYaxAhRCVkAYW9ffLGO45DxfnntVDghNf77NFUlcMQFce0atzM3WL5
sqgnT+oxubc2wgSOIdPs2B2q+5eQ5LCrxfete0or2RflX+ZErHk/bzEx++Er49Am6e3PkzKTg52i
Dbc3wFHl7SZFJDDGU5fcz11hX2DW58i2F95XHJ7ukC80GwApRMnhZ3AFq71TFVD9Nzp5GxtpHy4N
yc+/d2s56/xfIWpLgMLBZ0ILCpLmIvhNac7G2qwqnCSUmrSadRMvu/rY03fmdHVe5jPGZS+s8MBQ
xJlXzageWgcARukFqeSBfGfnQVOM1DDTRaY7bexD0bE2nGrtKH2z+maPuzM1DNXg4jNTaxfeT+RL
mXopJnMwhEKhIcgMcJ/HlVKayeA3+L6Nxomk1vPnQ9q+k2YXcfW8cz06JFvJ39aelSqr9P4c1OMx
l2wjYa6MhRtnFj7tNOK9x6XWM96N+sPdro8xbydAvmiC8Nw/BAk3oiTCec0fJtLeuUUdkPn2N95V
BMp0aGnTfTT0k22sI67I0JxHaaCHfjb2HBqAgBf+hxiJJUgC9Oi1zpIefIZP/07YbxHhHl0tRufv
A9/QJLehLU9+gaNdPtzigbizXq9Ze/TLbgXF1TilL6J5k9iWGCY/OSl5jqc0iUgpvt8XFCT6NJJV
OFDHU847VZMI5pYdzUECZ4Nlfkaw/as6zYHSmn3mw2ibqDfmjbZFZGDpqIB9Qsj8Ft+B7y89SPXi
Hd8kYAwy+P1l48JmQL3/Bc2hegzU3aceIYHpZ41TCqPQH/SB7jx+qIm5mbzZ+t2SbOvpvmEIRPlw
LTzaLHadoqDiNRdIjGXxGqNlUCgyI2cHoSHIQzUplVe+1Htdt4umFqNhUWDAcvc25V+6LGmhCWy3
OHbQ4e3FuctvLOJUprROJRLm/V5Q/q+nb23pnKF7UN5ReJHc3ew56e3hY7srZvO+vmjUvjE/8fmL
0lYaMUVzHiG10nb3AhbelYyXEPd15RV/91ZXpnUyhnmdauE27BLGLSbg+Ty13n0+iSsso/ZzBfdA
JdHeubaLq2BZemxZanjehc/jPOq5CJcU7+mYQNfcDmoH+V2lYiXzkojUBMWcDM2H08kze+Nq3064
MMWl8USLXcGtH9X1ksxWbdDg2APG5j9N6f7D1EcwjKWuStZw7N4CPSbO9Pl6EYvFRvq/qu4cCTP0
mm/7Y/iFINOv2Kgi5+W5kQYHBrmaXoylUK3KUzfZQth7vogZtYER587lZgF3VVL3LVgCS3zio0HW
rN5Dsynrtmon9JtY0N//UZvgqNu/y11WQ3n4nwiH+EA/a/JEFanwuML1p+/dfxfyCpYhTWUTyJCm
agUocbERjjWa24rpAHN6UJKko64ka2Tm82Q83JYcLcvRsCi/PjRd8+4VjFa8Hpr+XJBF6QMMmB/3
ss/Vgd0Qd6wfU11Tq5kxxMPt6cVMNbhsFJoFNKYUJ1ZI73eyOXMcz2JXLDhMEddK5CFzy3pG9DqR
DN2ND7L2oOvk6kN9chXRwVUzG3CMFGRnIAlmxCspOAxd0wLFcdPyi4rj92fafdYf9KMYKeP+9Uzk
AGidJToYpWUGEwE8BdK2Mfs35yXG2E9cg2R5wt07vp/ad0aBB4pOpnMzN9I3emiua/ebqccCnqyE
SgJX0qRjR5V0ui+FQTq+Te1OZJ/Lnk6pmsA3CNLZTpZya7rL8mB5kU8baByx5OzIgVlFljZsJntI
gJJsR5ez1m+iY0FYWv587AYo7zjPWK8GNL32puAUFpEWy6jqZCUpqgSM3tzRsYmzV0youjKUw+zI
TSwLH9I1pM3DBMg6cjoic+WuW5vcDztjbWMMCKBmNBsLFthEdsuvqYzN0m0Cw9B0xXn9cUQ18SVf
69+RYFU9lOQCHOTVFoYi5uNIxF+yusf6SyZ0jzGAHhp8IZa+n4Re6+Q+PQkbUbHoM5rmBoVtjIUH
G6qgz+yNLPkF/muPOcBa/uRPMciTFATmyXMIUpJf4HEOr31YvUSADwxg1aEM8CmSU02eLGvdCoh3
XcXoNdc0t3atdh0jtf6HIFDSwrGd4qiwdYFqGVXMeiiSFEc1Ki8blLS4wXSJGpsk7e/SwlxdC5ON
UcG4txex7+DN4uvOKmogKSRiPLNfbs+BTuC4i2v0W94C9VMDBxg//m2lP0CySSUwSWUR2Dj8g2pR
4y+NXs3qPggOwDrq47jtKubSduMt/dV9W76ZO3OD4L9/b9b+RSQVmAstdNWsaBaL3W3pLWkIUkX2
QNOZzrE8s9dHacKpviL7b5rku0a2AXZc9Jw6PS+1MjDXG/mWRxiGefxZuUDcS2mJ9YjZLxtknOPa
NdpIkU6pDuvA4C8HorSruVcc3OQBlTn8YXr4YaTFpmQdu/z8UywU/Vi6bSO/DrQ/sHicK+VY+u5h
XOeSdrRUYCF8QOz8B3sq5qFlU6EnkKSsIVIIqG2g0U96n+apqoLW81DYoUQG+P5tpA2KG3kA+Crn
u/SNoe6VQum/jsns60NiHQftBz048T+DIMgl3SxN3r6NhT5P2qhTjVBms5aUSoCSDoalczpXk27J
hoyy31r4Sxgs8ljZVtLqQSRJjMrFrBqnvhbNfhpWk5LhLWKe0yfzCbxcMifEk201M9YcfPDve2Vj
kCi03j1lr1ri0UcecT4t9p/hP6k0AgsHrP/7/K1vdzwSTd6qOMjIcSZo20xtEOxowfaq2OWO5flH
dsnRMTQ5S0oY2LDj96C1PBdYohW6snhwobhQje6zNfWO+ZfYkx2NSiqWSazIGBCalt3FOGOkHBsl
u58k1pevJn3/WyY9NAL8I736CdqxOfn7TLBGNg/TuJr5m6LkLeyOZRq8b0/UbJhMFaoq0i+WkEcn
Frtg0xEEqcU/152BomLnm8Mr8VoVHiCwZX44DZMVIlDouJYvyccbU4QgOVEVupCnNXP6j8jpE10y
pqJfkkjSx9VBlFobSo0Dz+ThZljFzxfJNWYZUU9xvWeyRyD2wXoMX1kGq3ruhUBSeKap5aXR04QN
8sdRQjOQW1+O/4OM0wo2DaniMnQ+xhQuR1Y5Rn3pkbKIGfOWvY3udLimaofZXSCekXuUtE9o3ufG
LxakvkrOXpWx7UPrISQjaPoqcIToOO9GHbGdRrN5Oi6hTiaz26U8KThn+cVw+NbEc3W+SYWc53vU
tFQczQ/fo2TKQrXiKqbtrCstU/V3E6Z6IRMhM3IhYmzOVtuUIi/mQj8ISGtvCRAX2WmMIyyjqdff
+k0pgAzuE7kjQpLJk1q5QbiOq7ID77uEbCGSlzAeVGU/u5OBF7BWDezgFyN09HyRLPJpBaFa+b2r
vCJlaj42CJekFhgtNYuPioRMuQlTqHt/H0BpGNiiNCasBgpUJEWzY7pof0MZO8TC3ha1qVzbfbCL
EqbOGGdwPACzwWQa0SuvsN8kMj2tm8NUEKXui2AiGKxTvDLYX3C0HB9ArjVg9UyPyrWNJ4kXNVEl
IfrslS34CXWhfrwnTD554pXcNBRyYwXtJUwnbXYpj7z/DJWk5Ahe4d6o+zSbFzPH+B5vzuGRB7zN
GdMQq3Jsiizv1AMsYlS2o4ug/N4Zxwflx1n6MxJn/odaBLttnL5Tpyb9Q3R+JipHfYof7SusEcHE
CAOmdCM7LVVF0spP5enYoICKDFt2Gvy2I9ksXj2KAZjyb5o7U6CzZv8X+lJRlkHsSK+jjcysrZB2
7EqsiI+38ZsKMgrXByoMkSqvZuffgR4fTtCLWrlM8gu+WOnnw0Grz1aeKEzF0kmPikU8YomCgccT
o2Oa8ImQXkX/tlLcaJy3nNqUNTLEnNvgQ7v1Haj9PkgZyyXMh3lsrzU+0U/8txptW17nuZudJoPn
nP5eM73Wsp4BaZRueqStVHT7xJo/cPSR+L6uQqJHuUdtlhdtEeLizXSgmuO4bj67b/pIh/sGt6Kh
K/cBz4yUXNoXmkh9Yrh2nFcNncwbK76lbVE0INYvy6x4PT/4Bu3msUHyrQyXHOr79Cq55LfH/1K6
zH3iKdCIeZaV81WM4HtnqcjIkHNIJlN3n1baklYV6phY6+DwpJeJBjr6xwqhoAu7IhLCuoG4Des3
NW897kH2a4eEidJb5FpZXvWG9p7ger+StfsCAmZiwQzvcVWTuW37vjhiVX4WKmBybmOer41jevJ1
Fb5KaA6TvslO92nVizNmwkb29GYzFdneHSecaW1Zs0zAeep0w5dwHDZR4ADm4KlVuRx0IyOYSu9M
jswtL7vJCUMR+fTrNc8l4j9UKJnPgIzwAcwFtcTItZppyrx8TjyzYvTIyJPncHtH1Bjx6IlNbiuf
jiZaTNkjt+/ecrZOoIBhhnjnkSvebn/aPPByOIJ+o4LN42F+eYEIHE36EZGkRL2okBJ6A2E3pYlF
l1aDdn/xyE5O5DCSs5y8xyEeDkjnVZz3gwD4EdQcgMpGdrBUti3O8yZXclHaZl1setbj/3gdNxVT
N5EYRbWhFbGrkFRBYcItBV/dXTG/noeZN4BAGHsQfi7fhWjDJt7lrIYIK6YqOLvneXTh4R0rSuiW
1KaqIOQYF2MlHa9SDMH9Y2ncMt8T2PYdtB1PVomDccEeW2+PUPux0/xeelGMd1wKynOTM6Ou6xfS
ySbMtXCvRujYsN4YjGO0OXbvNSmwPtaohcdpnFVKhNwIZluMjPnRcmDk7L54AAV5f/qGwDeBog0k
Ett0Ff/Ckuf76awHMR8BhO9iR/bQ7ZdNod3VSHw2cqyTlVX3H3BgB5WTEwsIbxQMBanhqzupxKmG
rX6dFpIbnCgUX5nF0xCBuNLY1i056cQ6hFhRNlee3sB2/o0M9UEJo4hESMM+qR1hzfG15E5d/25O
F4oKRqc36PGImKjS8A11DjqatQBsfAWtwlGFvKRTC6KcWWSeScG+/jZR0v/GPWnzVUH9s1P+A97m
VwU7AhnvvdUeG/Jbqg+p7kGOsohb0VGvlqipcMe8Q9mR75uHVLdH9zMs7j/Fd7crrnGrDnoTW2Hw
aLnZiW/nnYFxz9EUzMsfSjfVx9L+aP3JyfDQfoOC5mwxhydA3pYV8ROebc93X4Cflld/u9d9z6a1
17gbOtlXTXimJwEiCZLZ8gY+/omInNGC5u2fuFZqp8HQdLmbigqIysluJKFVTKwPAr05wxUMKi7b
eZScOI8OfXEwikxqoHHdQmF77vgMbVKupaTRcbyJMtrVJptIFdfxu+e0X2m3JSjzvF0uElImfTZ9
WxvumFzZjMHL6k75y1z/kfILodZtMPKiBDD/IHqmTuIWyuvHKaJqySUgaRjv0kSHvBtI1casOkBZ
H9qlya0p5dYaNhvbw9kiPnnFNLiQ7fhqWhvv+fsvhFYISoZ/r0GCSYcQDffZhKjlZtM8gJEtld+B
TSOVxjYHYVkYh7plfxdiEr8Y7d4p7+yNaWHQp3HClFJJs+D3byhyKj/BlO3RElcFikngoteDt0zR
W56gAgyerEUneBOUr7jEz8jGdctaNYMwl+Bcc9l1wZLPFQe79V8GWAp91ZaEQiCGs5XT4Ngkd1sa
ze2kQf8He0Q/QLWsPMxz/gpoCuny52WOE83mvAaVVU3cW+OGYeH0ul8uyA+/PEdS7zqqc3wTYuyx
rGj0v1b6zdKoxAEieaMgNBzpEXymm72KbofmST1o3A5Z3m2kYcgYrpO2kw5GJNSNWiLj0zTRhO5+
/7VAgURCKq4giSRlaM55wa5xAb4K2ugPAZ+YhHr7ehKj5zGci5JY/ZTKxVN5TG/x9rEu1a8Nob4A
AscQ6fSxk59a9tCcNxpayiEprD+Y77IxBntbLSIQbmEIouEn6Y498gYqsO7gNPnh5Z8A7giy9nyf
HdXhNstwzCdeLPxmWF996GSHvHoVyIOEhZwd0x+RiKxk8UVnJ/A1hltasv/CupB1ZNrjgK/Ry9uV
N5leam/SQKp3ACPQtSsmue2MDaOrxIxfhUO1iD2Uwdy1Seovi85/YKgepPKPGPi/y/ZVDpizv/e7
PFfNn9wlARrOPjYFx3F5kTEMnzBWna6RpLstsaxHc9VG2GIRttYM4Tmt+nhGoKCuj/tQxwF1u5KW
oCpidwFCQ0hPlpk9tQ+H+Dxo//gCBGtRUuYa3p8m89kHdTKdzeOLSvMC5Chncx78q0Avrvt2dphK
oCHQbEjVN+REbiSzet7ic9OsSjj8/kvFU/hOcy0mfHAv2iamXMHDpKhfia8UEiaOOgxHnkLTf7++
ktP0sFK75bct0/2WEw6bSh0Mmr5FX8JpNZsLR7fMBaGIlLQZ6T4eGTpXQ3IcqXHh5h/SLZ9ASCzy
U3PCttkVCDAebvlJCyVMb/ErvMv3a1jMBS0xms4u2HZhI33IfoTdL+cd5G5oGDzNsl1LkOXq6yZA
jbsnLUtvBbEZfbN3a+B/peDjee5crzGAnO+T2AjewlsGV56suwVdJ/wredjX0a7p2zZEmZ0+Jtq2
JBpM9bLZC51czKrLshM9cELKpnWxJ069E6k9rkmtn0adQs1F+VE2ligNCpUEbP5k4FlNfWt5it22
oj6lkpUWwDsEALYDib3g41IocgOws8K11K384VDeHtaTd2/cGII/H56qTyHNG2eVAcFWrIiGYZ+5
QRPqUV60sUjmGMU2+WPqgFr9RzlvmdtPcMIzoPZonWqPdFrdPQgGzQJ/9X9MEKyikRQWO52kasOs
1FvjaL+bazwbXSfoqdPoAVvsXk74/Y067PrrHI9phY51ud7899Q9GJpAnubdLtkHpzmuLBXEJlpx
enMZHWi6OpuOSZcY762iBb7pDnBPUuAtxpU743dG2hE5kLI6pUDJbJ+xkzOHCf/oI++ymGSRpar1
ucgqEcPGFPOXej8fCsY8TV0Yo86MzxgA5gSXJU6Xt1oUfv4Wsj9HquBol4w94ZO1K/3/QcJr82p6
QW1eivBjqjqzeXXDZKWL5AO++mSyTrQRNelTVIg0XKS4AQRldeAT53MLipgJ0lUpEDUmzM/kk4Kp
1KO7fmNo+NCTLR6quNrWqtoXhmrDGnYohZ8IObK0qtJDOFFzzCZKOA440D7rlJZBDKkHlCZ9IoOh
Z40Mt2guN58zrTrxYQHU8cYE5JS5Q1wAdFJSyb79UqgS27JM8eZggLe7RzZJ4Gy/W+9UEsHBx9Yf
Fd6DKNd9bhx+5OYnO+99iIsqZ5KX2ACXJbqojdm+Q37q7koHEsV31LS9r9alfSvSM1JKjUyfJ7Zn
vx02fHx9jHy83jELJuSYmRob/KYYJz/gfvawUDM6aO8AVbeRpkh0jSrZ8JybDs6lkiV8CtMAp9Rj
RxQvYB1LBodpASQu7VKhXNDtiZGvLnyUd9WPo4ETv+4NPXKtCtAvx9Na5XQohYt0AUCdAqj0uD+p
2MzLJJ4p6KrAUNGQLCwOep9281wcMMgClQMErG9s3aLWaBqz+a+zqy3I4Ro9++rTkRCYhzlKNDod
FoYzNI53Hxo/l1/HhaMzp5Vdo0vV9Jsxq9vLk8++R9o9PECIpXUd3G1pchgZRSy1sh6aVw3v/q7p
MxISVgyJpmI3DQ5Ez3ofkT/2RzAKuySef4OfjA85FLnjei1PUJ2MZ2/LJ+P8dbrg0PmqBp4UA8E4
7BlIEgTV5rrpxs2FrzbadFmY6MTx/i4Ohp6+rzlGWy98pwSGCybObPGOuFrU8NfEwbUa/yh0h7DL
TLmGreiOO4Sdd9KH2xrddnqjm6aeut/izixFhx+Flj+SRvbT/ImQr0V4GDBaFIcbJwEU0eAC/01L
dCv/njp9ImwQax6D4g/MMYm++gkrvJJzd+Ep8tA5mdRPtIKBCnqIuSPC6qeVjz8y4RIaIRIMsOW+
44GezFSR10Yj+4ya8CslHEnJNOEQQaC68IZAC57+t0c9ZT5vcAMfTNQk5Pdsa9LDzbIcNNquGJ+K
RhLBvoiuDUu5m/u2kc55JFqPu9ZWInrg9LFsO241G2H+hdD87vGHbH9kVHax3RPhz1n45v9C0bWd
RX4FKiFsC6+WhLFGIoiYDdJmZIKufAGwWOTickKMyTDxDsPjZVTRJdnReErmIAFgWIv6Y+OCS5d0
AmqAdmQ1DQ2nryFUBuOgFlkCLgjwjHeFAKp+aCR6fU3y2aZ5hTsqI83s8Xal4ZEtJrb4f6iDf40p
3ozacY1VwJNvbXCj6tHYTmuwxeWe8UVUOcD5zhOD0ms1XpkW2SE7yA2dTPCiKSEcK+w3O84PJbAG
9uYrjJ/wEh/GxwR/zKs/EPQWWPXp1eYaElopuJqafO4+6IaXPfESZZT66tCy+G3+e+7OKvV9hBFt
j3YAMjatkVLhAkV+czuuChkVLW9+8G7Ik5zJ/7DGcNwnaXELj+hu07CiLGX9Yy74YkPIDPsJgBpY
W96/2vqjZF1YYaR1rCRUunMqS74hHz5rpjXWLmSRUPHDGKgZruQawEjCijMexoJrRLPEyMNcZmbt
DeNE6uRnbNj/UH4n4ci8SOQumT0AkLTlyfYfqw6vBScIZYBhYAbV8pGYLDKArfDjfXDsSoY7KVDo
7YmnmJcGRC//nrwxK37Zg9hrz8JU5f1I5cker9PSF99OxRoyhtdkTd6sIR3npwqupgjtLur/xEfP
H8oGKWibG8k2D/KIaQakprhImqOR4rk2OFcFhG7m8IfoKiNZ4uFnqxPu2CJjxMWwHVQ3GaUQXJSF
Hy3WqHYXZ/MBrSoumOtgH1BOGdyGnIES5M9/WlpGEjNutJRkxH3833osGZY5orb6ES0rI6laDSXG
tj5SNpwRlTa0RVJCnt4Kc/negzTaUCPTvBfJrd9d+eUpR5CKfIcOkConSTHnFG6czSPNiWByAWGw
VZRUQsnIdgwjRfd+yszbSAxarF4ghbwJrEmGGBW2PObiI73YU7+XvErqRYlSll4cWeW/JAJJLw0Z
LcNRTH0W297B6AVOM4wbhbSou3zouLBtTsESkEazKlv+9j8z3+RQqxr3L9gYr4Oz2u9cVdFNA4d8
DYf+OBELs8qsJIYX/Jiz/xNFW1tLVrfFqtlQlu4Z5Re1/Bxh8YDdMzN1WiS+AB0spuehNSd/Y/JW
wW/CdyJ/2jOwP4BVJcTHb3ADi2otS0IOgbOTVly7BNFNHX0s62T6zd+uKSQkFyix59ExVUPCTOCe
jJ0TBXIpUcG4Ra9R4hdqKXjtW4mfPJJRhpjDtFLreM8YkNsRWdTcJX28umTyg/gEx/3dyrRRFO6r
zhl78gJl30C4ts58OHEd/IZnUGXytq66hur2Jll56jU2kJ/My0NpTUeZKQiW6YsfqnjN2UGrbvUj
nP4c1KNawnZpAPsqTwjxwkZ7eZ6yKmp6XFQ9u4Tw5Vcd6dFnGxMUG3U+JwWdgB1MIm5vRbLtKc0a
XEJJxOtP3FiJkb4EdpUDz+NeZvWYX8l6vxQ5QeHwyMf2dc2U0JtfV9zD6ksi5wfL6UeXt9tYaaQF
IpK31tbOI8SUkzSPCosNvptXq2i5LCkRXQf7TRKetBv7Od52j/hfI0imUAXVPMBjAb+Pyruwo94j
4aUIa7n/xnCLw15xMpd0gOJ8BovlzVTC9ifK1t5qnQkzIdR9uOh7m4ojIPekhfC8sXVQRB80xrM3
NEOKlFe5uxGic4KMPxXSRtLvPR+uS2F/2wLaqqg5nfZpBV2JyaWStC87sZ/JS/TiZ1zxUvX4Sg/n
QUGpwQL+9iH5B0aDUumFq/645ABewgUt6eNjw1YFi7UFAOfj6vVN/YVLsRRsqUlj6/g9etC6u15Q
kT4ktnu+EfrDLqpLZTnRUKzm0EvLNgDbapOW/fUNCVvyw778toJZuXTI6xogQVBoaUidsqdi4TWd
mzvjoJ/dCPtvdoRTUPHNq5wOYlLntSYPbQCTiyq2T8fp7HFVQ469tTqIvvGzVwTBM8RFRf6aORQF
Hi3AwoLGHRTeNfsxTAQ4No1zo1l9zs5Go/+xnmsBpiX08LyrMvSCkj6507zR4wS2xHoEELKtPpDB
uoZmTZSy2ddV6KZG4uWcHMj6QcYGce56nZoZWH9YjZj+IwTrEa637tYmq/z0Jq2xO16ssWQudG3r
TvnFG09U0Rd1wCPmZfMHDX+keYAACxboQD3pIElCmvOmyC4wGoDchCA79z8vk4fgf4WVNFUautLa
UbwMmlNotl41eEQ50rgOrYWGnW7P6nYtwubfawHfKHA9ckAYEcjXJprBXBVSCke9VaeWuB1c5fuU
QPinmzJ/7XLKhvdwrFm1jZ1Gm/lChEAFfbFcjDkEfNfSMsELaXdzA3nuyVyvYOosWmHMIsMNUhim
rSrkERBvModcWkxSIxKMO22NcSX9Q6bYjmeeWSuy4pLL8L54oKEPbwKPGUSpX8hAFHkjXK3iadS6
YVN012G0NVcCGP1Wb7xlBChUrUIVfhuZ4R4CHKcETOuMLkdZofRApDcRwQIP/Ufczg4OOEwS6GOm
/L4UCimtK54/2RpizAvVGaBvUaKlYBXuyVUUwI7qQ+FO5gIVD/9ybgpEKdE6o7zrz6zpxpHe///L
8azRgZnf/uaiW/YcNR4AvNogSTr8N1uYL9BADp48wxilBday5HXBDeFN1w8yTNEPHINZlmYiGaWx
SfCT8Js0XzdbO70eDvu58e5RJu/PQeP9elRt5oNBwNP0NCo7qfXRAPnSXbYz2DacteJaTSGThpl+
wMl43879cwqxJsbcuVcSD3l+9Ek9Q7/u8HDxAY8c75GDldapGIamUTcspvCxEZciZko2kzbQ9Mub
PgIAcxrMtVyWOiEDmuFyEYdYdUZtQo7vBE3YJsSQf33fEwPlXqcsMa/aVlKMk8X4atCv+ur0KhMy
5t5HRFytOE98z3aKeYn7vRzKmPXK+tGWobQ6MMvKOrcaVAgVkdpKBxomqclpB1n5nGxIWLgppFRl
FaTyq2nxih8C+O3Sq+a1vDZrFj6g1XCwOTdLDKgc+paBmy8lASEq+Jt678XIS6za2OMMeqBmT6/w
kIZKSmaVosAHAZcaZLHi31WA5ikUA906LcVLw2MaaepdO8WgcCbsPfmd/zeBWO4CeYE8L6tN3+9A
q1/RpnO4DS7F3c6bqqKe9sJca//IAldJCCEySZ+8pWUNieTdQtG7LpwfnDnrJGjdmZIYB9+8EZQP
4IIajtnzo87zNdvmKKR0Z/lkt+IudFm4J+/iWgq4Ya16e/Kw4kgiTLTqUy1k2V69DmU9uikqBYCq
a5ss4SXT+DYXJLp1uxgzdRvb+iKOgFnkhGN7nWVUd39o2GfZLqiEg+qwjQkNa62D+tJkr2xVDJPe
uuD+5MiRQs4umCbH0ewHTcbQTj4T8ZAXsXF57gPzDB8lI1KcUhGzOKE9eIF8yyU4fUMv2iTiakuh
mBbokpnEfy66V+0qc7OmfLlrJnE24Fv6DBmA8wh2emJ1O45gMGgC2zatyZsajHT+l5O/TMAGfe67
4dvvNf40RTzN7JCVF2AJS0fQpQfgexWu7FXkiWeP5D1PqV+FzfZ4M3e5HFGnWqPQBFecQh30wplF
aPLLEczjYiGa8guvJRjz64NCFPS7HsrZuszWLTchqtGpJP+H+3/AfKnC1GoPErQpeBc8PL40PhuK
NoyEJSfUs32ZIlbxPlmRh9EvZvuj1o7V9Wy01GVbo00Op/psougvEyb+sdJQ2u91dA+dp2BZr5BI
X7EZZ9+r4lQzdqVipNaDsVgWC0eFps4Hd8Ad4GC2KZmYSlCEGP5XRB0/mmTi1B+yVS/bwlPNGREh
74a8sNzC81Dj0QYqhRRMOgQ+Z/wsM/7juls5qLLynmx7+YnZAMqRrIFrdLH3UQj0Lfi1Yolgm+ny
aoDwx7P5i+buzdxbGUVtnj/BNK20P5QAOXOUWa1JtPytdvf9tA1tk8vQEQpMlTszUq56/LniJyZ8
W9aA3fg2i76J0ygs/1HlTnpZgUiYIl2wq42OT2qRINHMt+jHWV59Pn/iBe6aa+AJ6SuWlmiicK6Y
YMvKmcn0Io6KoEayLy0SeqwvwaaJxbglhhtqPVWPoKR/fs/W318NwSuEmzO+xbGAN9HE8Zk8TorE
vQzRKS5FQBv8/xeO4aKcng1VEPZhBSnVOXf0YqXl2fbUuVndhbVOTct1jVO3HrrxQscVGTjCgvu7
IgbTX6fEVzJffJujkCz5zxbmXPfmQcg6aWlO+YH28L3GvIS74cc1e//SDiLx6DqL80dwmRaAPrKh
HAbSUDfaXdhkcfsAaC2t7SUI+UWnmKx8tqTTgKDkTs8MmczOclzWRNAigWy7EZALMzGHDnwzXs43
Gwihjwlndf8IbFS8GXI4IJsuw9hZ8Y1uYDgh6/F3le/VKhv2RABThjHUdnJ4pPjhYz2/amjOFFwM
yqsKYxQ6a7vXcKjn9j1kKDtlteqEwCi/zk1nnu4KLB4IvI/2YwMabJ8qDTnPM3JLIoJm0EMN8HJE
5WKpQLSzw8HGF/QtKQGIKBMElK7snlujzd0JuRBKCZdlP2rgq6QkRoOMrUhhmRw/Jwyr+JuPqi3+
NuBXgSmj8Lhrk+SzL8H6JXMfhdQJDV/vmA5uDConjhwzPW63bM9sofj/e2U2crwcW8s+xE7+cYqY
78LSVJD4fsTyA+6+oCgChv/AH3eZW4a07xt+pu3sQbUguXPG9rxcEZJkI5voIzT7bCQseppqrcRX
YrDo7KJtcJShz3tfBiK1gryXq4uO4lvCRG1PWrGlTZkAusUb7oHDVCESDxpLJCN795sfdNgxxbc5
5jUHf5dRnLxA3qLokKWVSs/2EI+QEGl/BRskD66nywCxgH4rupxTeLfyCQw734XgS1JFoL0x/Gfb
jt6YWlaRtoubZLNBn840+zRg6y9Ay9djYrQn9XcmORJnFJQk+0/V+eKvI/9P58DAdzUWckVkzcvD
gjwBmnEwH42mx1iHSKf93BsRn24fJbmW/miXQsn5NKQNF92Fbpk12oOir3WT6cdXKCh+WAjOXk/l
uR6mNB5EoS1P9rBgIvAgK9rR2XRmok0e5KQH8oZXLZdBSvvGWdhcOljN5dT46YRAFsqnnCf/kNoZ
g/bwqcyDPT5kTDodey0AJNRxE2Wy9qHWaLLGF+3WmmtEaCi0DlS5UHaklmDkw67XUzvq/IyM27Gi
S1q0q1JlV/t4q3mIyLrCixkA+szipWUCnLop6kKGr96EN4qVCiNYMgI6jmkoZdQxvNHowDKq/YT8
2bxfUosEfVBIGdUGAnewuc/+ApYE6UVbejQnVhCRdaweu1sMat90RDm6szPgrlXbQb+k4/LMm+2b
HHiSy8BthoWWManPRZoaxmDk7PIPgX0Prxg3H7H9QZBCDcKfp/fVch0dX5SCdo/wrO2GT+xzuiVV
sI6u2ctdHF8JTyhlZC0685roEyPxhiBHlZ0JZdOe4QvvfWwi9fFR4AkJNuufhK9FfYoatkS0LG0d
rV+ZJcdgutGqWtDs43nn3D9KNLf1NSimy+daJvVPhGXVE35tas27ptMNBV+aaOtzY6f2lEXZW8Ap
1bqEQHm9a03Rihf8x96pSmG1ssby1aqkkIwjDkHemQsUXuqTRZGfh2D4EzlVTbDl+0aprWT2cPeR
Uj7CbXdLtRhhtSJBDrc2CtM+QUXDebzbmx09yS6KZbjYOD8BpZFRH96esA6u9XQQZ/J4wNUSXgHK
rg8Z0J0qO5ICF1ZDj4zFV4w7hor2qxnnyc7oaV+T/smLmUyrdb9ewO5lu8kOwykAvMxoIIG7+uGZ
x5AMFRa8L3V/qYUoxvwip0rMgLg7lWwjniCsy9SdT03ycYB+WPDm8Q1yT8Vk9hOpcOY15hchB25L
V1+drC6JUDV7SHq31k4sV344BpRV9KlNYJom6HMky/t6R135XyTh1b4aNKqduK4Ani8brLT0B1xF
n4+lI+VDVTojQlwjtNCzY4ydKhOaRt8zYwOiLR8wDsYeiuXbM/N2eA26n1yOpPBQK6gAcb6Ti73x
uLUPoHxnKTMP72mkcbnHiZkG7R73x/jAlmcd0XIc+0boIDCfvQURZeXTuMAH7qvMKVxRPOoc73Ms
Wzg3BoqKj+5lH734L+cICoj/55v7yLvxSV0gEF1SIhQGUaPuvdp3Fm5x/A74zhExz1W5k4zdBLn2
S8pP0oB8/1tzvmf1L9MTeikb2OOxxQ2Kod+jA+s4IK8pP0GA6WOw0wKCFMHkCIKiQz46Hocn+a7N
MoXi7GflCrvNdlqaj26pHhEBL6KwUNOL94vEUJYa5l9Js14PPioeojT97+nXD2Keakb8/Kymem6W
AlzN4YPocOS+oU5NKYhznlQWrWaPXgIAfUCy71XLJRbGPblhvTgwmhPeZ9WHATwjKe6FMVOOUzrV
HGH86ZLEkwXEWXB7WEOtc8JxqEoN3u0TmGkDrmZpGl9vYe/HiSoo/6kYZq6tb1dwW8X0lFLkTlnq
hw/sHCSg++J6Le9a8eHJgzxDvcUROm4z2ms33R1VFgOp7ytvLNRcJfqSpHHxCMd3N2EtuLqT2Ggy
VNBnBKEudU5qQXZ3XQexWxGOmQQesWhsXOUIeZf/A013vnbaPy7h3aat6ODUSE/rQbwVMp48xJ69
Vcqg3gORwtr/xyHcy6x01m93mB0/JIDuF+y8H/dH8HqwEoNRIG22p2IaWtsSN8zxRUrq7m0IOfJC
R+0/5WSKcQhtvaQhZ91xsjAyQ6ecJgQPYAr/hM750v7tID1PmNrqpHqBASSvfKWXXYpvlca45yyZ
1OElqkcC40QpZhtnoAgIxWXqmjeLyCMAChcMTEwez+T0JXLpr+F73QV5sO4SqPJYaeeDA7KhrRBa
A20q1ct5bfYKHbTMYzZtGE6DVixmq330KDpqV/JBxuGkxX/LdrV2FwlPIh3HixSRUu9gdtvPiXtv
6ZVrYnuLPV3eelQGWzk3iTgKszDItipn9t1VXnqJ4Q3CPAKW0BP+RGJg89rxIv4GNMp6GCwBEalG
l9QqI9wS/11tRDwkrovhsgNPsiOZ9eCUaS+USs6JmFn/WJbeBPYT/DqWbcUA8MJxLX6C5DHlZYd3
qf+pPaMif5VOiqVSLFR1oawZz/mlahQMDWazUXfe/tZ1xkADtBOtRmAGT56zsRN9+MZCqtsCSfqu
N9EEYIaYms7mhoZ1DOPCy56XYtCNICl2RnClV/z+f+/EorVPFLwmJL6Tp+R3SjRr25+yQWPE7U5i
kmIwm6dDhDCWnNTQF4G4reevmClU8yuagOtjqjdGOk8MH9p3OL28+DkvP8OYhQZ3ePfBAB8N4GeN
THqA1fnbzhZF6KSQ98rNIdCACXsyTuuyk+0vN0QZuIVlgVwGLphSNbBFVqspeFzphBUiq0+RA4eJ
ig8kyFQgmYI45h54G+tKpd+x3loA2uXU72/MQR12oVdeim7S/X9AYMNVnmtiZIPhUdygC85YzzCA
6OQCSkLKldQh0UoqMCuhbKGKfWWGn4sURHjVsVpsx86a2UKITE2R962lJMzC9u2DBpF+GDw0ewiO
/9qoK5H6fIH6YEFFrdD63TzRzPrlgzl6CvKrPJc7x75lw29rB9aaOMrTIjenhvPCOeQYTiuMb1UU
i3rAGdqxMTt9L21orujJTjwYUrcAyXgVDkETmvHOawwIfwuIgFP/W2mUdoLn9DB1zYRl6eyqdd6K
YYB2moCLC6AgBH2/tMcw+U2iWUP+W4sTJx+Rf1kbeBZpjZGESzIZf8kb5V+cbdyZa8KSMDBRpVXE
2xz0HqC9gUJoaPbMvbUliqob+GdPk0M7izbWfptuNxEXuHrlth+Fau2+Wu2/idrtnB77fyLquw0X
JtjgvwUNE9DxXY02puHw1LlmD0k21VfpsmebhMjulrQzqmByZafI09TO/E6PP5Dr83YomGRlNI+Q
VH753XiqNAc4PUIQSVDaoEQY8yuLXNov7CfLcnYS+Vyb5jOZUxmzwOIyqvA8GM3nmz7Pee1cAs1C
qSezzmClOdPUjGYmeVftDDP0L5QwQZVXZ5EONo8Vz1xOZR2DivMo+b4Dt51BB0YKH9MCT9Yuxkos
qc78eTDfNnecStGzSI3ZAvYxVyKMATfSnH3f6gRkpN8HUobvMI4ewrQil+UvUlfqR2AbQzpxMafy
9B5Bzh9ygvmOb1g54Yz4msnuStJVLQsM8M+ZKBXUSiwM1XAx3u0D8PuxrUvRBi8B9oVaM+5kUnSb
XfjNe+Z4aVuOQJtvC9LHh0TLsRXkmRW6Irb+uSgD9flc8bl/GG4Rxd0lfzQJMpE1cq6yYGSZ3se/
kTvPXiohlfarxIvkCVvI54zO/0fR0qFd47aAS0n3vKpK3sRqIVZ7p3BBpftYXO/jhYN6FSMvGXUy
DOLt/IC3ZoH8SAuIdWoXAACXh56IWPDIzUHfh1rqeSA7mwQBJWdl+21C6CkoEZ3QAkDY5/iVmsSF
X09pl6Cvdr/RpVLbvmqqi1hO1uSppvPO1lsR5Nri9L2uQwavYAy6AWIb5IXfMDjgxKqfDwMF3cND
9wf9cTHN/s0z4EmMTYIEDGqPXIKnRSr1zhQOcVBV3H4n8xpTIDJ5ncAa4n3MkaK+qsfzRrujhIP4
cCzruccVPFPx9IIEZFS6q5yMLmmhhzMWViWGXhbvQLGymnEx2pK2cHXLdab8pGh1j7FR0ejdtZG2
25aMPIo9pdfBv6r+aXerFZ7qZk006iZji+SRZoNVKfNrQo7f7aRFuhZ5mJR8YSnx8vr0DYocJgoD
KgABDeoKXSqOz6vFXNXrgQfDPGEwx6Hg7NEKJWuJ8ykhfn0DmwICBdevXhxL8WBjqsvr9DGR20FN
1TapicqYOaxfZBQziwA+UnTnePrAiOidhaFl0Q//Jjsu5vmZnIFu7tndbQIyb8YZ0IG1Fe57S0y0
aPxaMUmnyPG/ki5zqZM7u47n5GjVMmdf+YkJF7vds8FUPXFOa9k1v0MXhAmuXu7L98uUoeVt1Da7
0MlY3o7pVFK22mo0Mis2fguuJtEyIDySwFLbj2kNbTpwrhS6Ot+ZFk/5cCyAwYIIA7KET8km9vMg
UTmgEDO2LjkimoVu+0WXh+jU8MLdIlq6sRGDiVXnk6KnL1QsdtP/iuahP6bys+wweymiZeXOt6bj
6tbWUDJCz83jjDdA7jPJyFaG63x/H3VWD+Z0YZ6G3XKtB2Aw5kLsmlSGC7Z2i4SIHF53MjOEL2YF
h3wx02WckkQVfSHa5QKYlYIGEgRns8tIvZz/XGyuE8jhk5xx3UQEkHCRP1Ue3eHqYkvUw9jy4KPz
HA7xtTLxwxjGJNw1WEIHhyWFEUEqmbb9nQh1B8unu6Sxu80bfo4MxnL4Wu1M8XHUVJivi+b2Ybxc
pxgE11g60EJI9iO3G8uffqcDGCCR3nlduwHk9MI8qmQE2sQQ0KGrTqa9Lmci1YPupEjZ9mw52sC9
xHCZkGaNPjr+tHBmUKe6i71i5jWznKACwcaF+6u/eFtzJZ4IFkxn5/G/Kl2QjntThAYp248tXhQL
spNzsGemgEoMqwPrSQICKIalsg2dSkYHEbKIQgiUrff7KG8zDSjb9RKRJyrg4unLh9HmYDSnqBLn
FbIJ0ZETRhYjVyvNrLoI/673hiU/0ZPsa0zzFPe4LeMXbsnaQzpNfrg2YDBebI34uOJYisUlgSyy
q2XZqQ4Z/gmPQTaLv2p4zSuwOuLCZ/MH/dPyCXeeZGgqqVwcOSxCLvSmo3vNTPz8T31P9Dz6YnX7
2Lsl0TXWofJcwTNWiWDEdiAAvwpdWJnMzoTe34L43HvDDUKH/N2cS1V7ujVVsfB84jh2XR0UnnrW
JbbVcEmY3gzq0Y/2pquc3BwTBfIzTkGnokCiSaZU7uqoVKy8EVQjw4kA6sPaM8A40pcFUIHvRAqk
K+uS7WPNI7EerwJI8Joxmpw+5P4s9kZTSw9sDaO+kJfCWA3p9BFLMix00UuvlfofTaFYyMSjBtfO
4qR/tE3z6O/oLU53ue3or7Z64FVoQD6Xdc0IMWLm3bb1ZRngosz92VTSJGcUE8i3UUlJncFuEGU3
h6XX/8i+uAtZL1MYiOXJi2yhOaMPWDbVUr72c8p7g6sjNC3FkpAcHcw2IVD+3g3pBYdJ1zXD4O4p
6mHbKy+/2bqLmWqJCJ9iutnPGla1vHcPxi7n254GuXkxZZJHn+kYLZQ85BK1+SUCOX2EnZrSv+nB
4T8CCpfgt5pVyyTuFOqc7fQqcfomtPx5aEFDwnSLwFRnxV8+3QIqeSMAl5u2bIhgdoeh0loqWihJ
YTxIVflXxIEKzN/SXweZzTE/5xXcd/8FKC1KRvBZOoTU1Z4KE9i7uA49iKJq2tI2fFe8kKHXtygE
PorOe501Rnu0bNJHVutwfznspvLTMf55FeG7RRGdQKCZBY/QrJWuBHV8I3SwI7NvVNqMENA3tr6Q
uDwhAVnqfkZuE4NEIAtc5qk18FNFdTtO05XE3qieRzzH/LkkByuEo3VrdQBblGyJej5tctYVc7y9
hLiL7EiDQR0OFVRV/YhjLYzMmgzlANutNi5j1SEKNgL9gJqfrmfwmVSwhIJ2O3JSM0dWai9fmjjc
8r/GSWjJohh0QMA+wHyw6Xgv6lMPNjMJa/j9J6J0FhWALbFo/mbPGyoxJqKnb9x2sYkmSw5XwNt2
dUp6kkWuQYe1nTjzvLaJLMoeXSY7icu0SAfHrtRgD93roIGzxZNCpFxpG76TRrlkE3xhDk/gdF2E
58L9Oq+H2NIoENQx2EkjYF9tCnxS4ppuWgs6SjHbfoneoxvpe1itxa1dvContAFObGnv7jW8HCYw
zlsQNVueSsQ55po/uEo2WMn/17jcleUJH+7e5mUjW1BwBID0SDd8ag1H4PxiLj9aLIOxWuth2NzS
3P1MZntsswmONZeYBqL7VIQ9AM8Zpi4n5EtuRDaDwJ8Zcyt2KjihRKaUc70kjvdyT3JXjgS97Eym
wIzlqpZU7DL9TAZY3yP5UtPFNSyiWFTHSaMcsEwgkUxXQjPKFN+GRpMEr4vuCfFOUXPPLS9CT6yu
eRS5KbSYG4qoujD+qG1Ajj9pJ4/646B49BO2/BdHR67A0ucvrJ0mDUYciw1aI85+8pvdKCWce1Lo
l13cvIxi7dJDKrQhpwfWPpajHCwgoZNuhWnOgNY56htUcTqMUEitku5rq1uDdxBwDTf2z90hlO5L
puQ6nQ0XDd9uiZpUbvEfARxOnoIE5zqXkHx+ZZjexC7UlfelOTdNx3gYxAD35Xax5APzSguNdZ9o
bb81kbjbp8ZS6lEkhAyGlDmXh6Jb4l1NCw39wizdWFYHbSSoAFzKNvvDp1hiSJSCtBLc81KvU7nt
5OgWF3dEf2M07it2TaPTv84ZE360R6DsTskv0BI2tvIU52L2japroR8U4VgTfAkQ471UabQa9ibW
hM5+xxgfQFXR3VLEyJkiEixhIa0fQqjnYeedWVToWx9AXFqwfiSWTBmR8SihValiMqYuSCMbG49B
CYYqmSvbEGrzHqcXsUVJQDDLJlzctGIzIKTmXOYvZxt52GXY4zj5NlbtFUmIK8vsKJybdXD/WA6j
yqqAW81uunh3K14aUhfGpdOtljZv7x6cAU6SdY3qvolXI2YQRZfb+Fab6nnSlJF8mfKkRM3Et9d/
mKXCXnI56dzvIsjC+TB5mJ3fEzbXRAEhsx692rfunOEKmQWp7iOZXfkF/NqDJvldjhXCZvQtbKng
jOjL3dz0du6T9HZWcJwlqUcBe/6x4X65rIDwNbfe2GXW9ZciV/D8B9ySEntKVAyQR9QyxEaHySnk
YDreDTAXYJJtBWtzsaW6XVrvI43Rjwp4/n5X8ypfxZ7P97dQH/GlvS/Q++qBK6dW5n1qtkl+KEdQ
Jwzuep089MPFmw/+tB7bBDyPdWEELk94hssjpsZP2TJ0YKMRZSXzc4KryTm/jYWzKpP8Q5ZAiRp9
gwGHz8WyQZ0CkQ4s1JX8X/gIuVfAtFgaUGlBzIQBdhLEPNDGCyHxGx34rdo9oYkmlrGj8Iz6VP/O
JHbp4RssUlFV87HJfHp9dTDtNPm+0kFj3ScT1tbeGzarbAR9gQEP+SFkwIDKJCYwXJWv4ELT76qG
oxEJcuoSMdvKzOTtU1ulrr0DAiPCe0y1Afl14vtljSUHjvmVYpb3LESCWR0gO8FtdFCFndUFrCKW
hIUsKaj1VuY2yjgQfE9Hrv5Vjm7kmpDzWNT9bvPeh8suxlcJJJXvxtcVxrcf6EdBy4oKmeWxZCyZ
+e//dlyC5yI5F7S85BIp787E+OkX7TbZ2GL7VePfpODjZG6af8YUlN+W1RkgCr95FrTxV2lMi1hc
BZL4MEdxWO7Y06uEDSd3BGETMJ1sl8HzLE7mGai8CvLuDyKdBqGLVeN23ezGkWj21aBYQgKY0eAX
g9Pi6vn1KWRFskcg39ox9UVEFQcmd8Q8QmW+voVQ/2AftJ/fEz8SxFgBwD7PFiEzp0LQjduM0JZT
uDYIOaRsazgS9TmHu1XHhPmGB13wV1tieceERVWheiUxxJbW22DrkKdZRecT9psn0TyzWVv+Lkdw
HjlpPttsE4s+gBI09QMd/79LFMHBvEU9S3Nh9nYHu5spjJWmXu7mJ3xhWr1r4nRzU1BNTkgCi9f4
BLNj0Z5rxgzaxQQATZrqanf9KBmslL9a6tLRlq5ToyawuFfGYzT9mW5+UUnQh2dACpO3e4lKIqHc
FwWDPLVa0AHltlfxoTFBcJF023MhAbbXrpXcIECe8sE1bX9UrZk9qCW634ycW3ylLGPZynhm2tCI
W7/aik8cRxk2/0PWfNXbmEbLgN/sMTZnkxm4dfKZxXPhqPcR5m7QFOUZ8UHWBZR9MhayEuYxAss8
9SIjrFXBgrjuUpVYKIuMMbsQK3zcGrP0oiLl0ar7A/a7VTjk7LRzul0tseVJAViasdt4Tl5iHcyt
O170o480ETErukwYl97zNydSAcBJk7T5+Xz5XXdaDFTFLn4wfeAj3CFGhnxUNneBelLTiZl3CpnK
Lcw+RvGcLTWRGHb5P3QQL0dc/zx8Fg3tGVpcavch1Gfw1r5oaTRKMOt/CZgid3K7V4q5fk3dcV5j
pvU66+StdOZgHJntATM4bIeaFxPEvUzFXN+Yhqs4eqBOifNvkSDo+RKQKj8b3QTNNNfKc4r124e4
Oq04gcRRmyNd6dnbo5SFGEjxCYrCVBREi6tKC3IC6YUAy+iU7wSEBpjWF0+/jO5boS7QVUwSnoCA
37A+0wPmhipeGwwvtuid7Vtui/SN7QZuV4LewKkOUGnbGb/ZCuIglHvpmp3wCt/3LEsALuxn+jfK
4JOUhuOJCdx57QWjOeh+eTT0e+J9yxIFqer8WAGMPkI6FAT359ZXmYx4rhXSGXsVPcwyXVOVTsO2
i2cIq3H8jMDbuQHmIqp0dOqaBxzc2pU78bb5E6S3VxomS/8te+hoJKWRaREH3NJ0TOnrnmdPFq2R
rUCKMqnoe39BqlWVS7H2A0pMP9XXq9fHpA48ZZSyrmUKqmFb6CVRnL01U0IFz/0YBcYps89H8ndE
c2u4+cW0QCRaRqvEsKPIApbBeM8w3X9WzNOciFpYGHJyOuQHkeeTw/988viczhqOtzuV6TR1enot
EC15Y8RSIHXh3Nyyg88YCGAgV8LWg4FP3enEPAu+yARKYhl1eg7Aptc6inVgZuZVIJU4XBV5WRbJ
suo9FGGkNKBc1X/U+PpYQOWr+R9NjGv0DNm43GY+CmjJmyjXiGFo7/w9dn+QkDwjKSONRNXNKRvT
0JAFbcS9ZRnHDH3OSBaItS1CeBcL6O6s0lHrvwj8zNnY8f2DbVaN9SEInbem79KWcSJ/G/yNrqMD
n8PMOLn3ADXUTuLg5JFV8I4p9WSmhw/VAFY77pQtK0QsTy6ElXelzmw93+rTgBcTlobvktXD7RgO
lAWnfmcNKQ0ZkzwwDS4/mbWit89+vuc0M+jlnfAPYakNOaEFmQx4zMyIYzdo1OPVhltAGQkUakOU
9a7YHrkYrsSj0a/PlArtRMUpv2xKYZWX9pbiYU/gmOoNw/G+ESd/becr9fJZ2etaGQ2Bm2KmCoNz
nHgueElz7P0X1KB3Hu2T0T59BNVR4yOXnJVz9jt62RuuAYraKGN6dLheW96n4RkFlkO5JvD3sYkC
ZWz535Lnfi51NuLKFpsEDnsdgczCJPZizduXoH+5ArkiZYfljPPweJCiY+LWbWZFCXWxxAf/OHna
adwbDArZmPCxVWWxuiZx1GmifpCmbjuOqIwTDcuXG57a2t/v54I5AMMdMkNRTYyj8KyvYW/ddRSZ
7m8cMqmug1HP617yGzSXISF8U3uuqKgfY8HzXRIQz/t6CucWIyVv1ZOA+Ccouni3c7XxdbDDetbi
A+lNBds74LH75Qjcw0a0GCfiHwXkbLVKPZyEV84OIqe2YE/Q0KFMK4Lbny+hGHW5f1peEZ7flxfi
EZvCn9LdIuhDy5A1bygs1L7pQ9HzCe+XI2LtRZyPiB1weYek3siT9wQDGlB2KehmCKaAri7P8P20
TOq/Wk959TpHYUwE/TI3QO3t5DfsXZeMy7f4aDDliXjot4t3lR8mPOSPa/43rujQvLhGwEiQqHI+
oaLYyhEHnK/KRC9rbCxSbwIHoFAeoz7rSaU9n/8tOyvKednjn0IK+ndhIxju27pRj9wa6RR63c8j
2tsfyUUVSCzl4rWYdPk/nlwYQhT8V9no9atYCH0/l7b7khCyb2x0hVSZ2wUqAdBhbK0JW/Fgu6IP
kdrXwVo+fMqMAc4IxVjnKzv+hBRuWXsJvHPTkTNd3I8lDf1xxkEcwRMdp8bkGAVhgAGWwtZTSXXt
44fParoda7uPY4EOsusxUJiQhwfDUyj1yq7iYnPBcA0UumjFc2LaHv2H4NgLjQfTE4yo7IqZCVPM
speQWKzewEX8Sf358Gm28Agl+CjHMu+TWMaezNfTUnliFcHeWPVyyZf0hYXFVyig4ITMRS58zqWQ
vJWj6oi6/S6CwN4Ydlph5nirR0uZM1HikIa8mVDPod66dHzytzq0gGHJnCzvs4mwbFz/v/Sapu3w
zGRdkjBTWF6zlbtWFWvl08azq+EA5qUIf5Z0rh0OBcZNJHHx39SOLt7ijXpoOXv/VJuBuaSIS1BT
6bV9kQVNSYg8Hn0Jz8RcTujAkVGgZvQIp5j5L3ECXNP/qEM3nnaJfgRVy1PG6pXDJxAUyqmcZKJe
BlwnFb4Q8BDOaTdfUTwN5WOwoLn4t/R45+/mqfNPHUraXE00dq39nzgFXSuUdjisri9nizDwW5t5
w9VpN0Y3Zu1kq36pXcHFUS/oVtMtn3wPJeUpqzmmrZxLfKmQ3cliwbYPNmaJjHerPHL5ZrQPh67l
nQvTqnB+MrATs1EBiNC7v/2RaVdk0ZixfAqaiWVkFN/HyqUGD1wlNbwn3mtTbPbxRPYRwPg2944A
2b5bXKKSfRNJZ730A/EkigOPdAkkRJZwhx70B0G/MH6hk7WRN3LmhsC90o9e3XVNfq2bvnZC6fNQ
xs+G58ZySqMAiLINdY8/nuNLRTddAPWuWbRSQ5V5fFHzODXcgCear6uKkdqVMRo1llbMT3PigYKf
1D8ft2mqPFsDyXHSn+Tf4fwGduNnUI5PERUFRu0I0q6Nu5JNl+KV2/iaiz6gKHSFOm8080xznOV/
68/ZkRdW1keohZ7ou0NrDKY6chyv9ufyX/BKALX5I1g5hX3fQpAzPDk24mH1hxJLxkynt5PwuB51
JdbsKAJp5Iw++L3/hEljBj3TEuTZ5wKua1xtIrSCFsNfLSpvUBDooEItOoKqiigw9aUasmKmQiOD
+SwZ+cMwUUcGOcWA1NWXtigJWaRkhtD+Gtd0aMqiC8Ky3h9kmgv4oOeOurEMI8L4N4xaDIy/fzAj
liWy9blKEZNVu7VvWa3ayYoImhVCvDOpDWjjdVJBm1R0K9GT/KjptbqbsWhUJHPQvL6tHEQz0Z75
RmaTeW3ZCTkvzOIsHQM8kpUNFWXtJ9ZPBdS3ObLt0cyJt9QLz7SukQiRRWSBTp/F/tnx61SQog/q
vHMwcG0rUxpwGFJBlF40VLVT0OSjBvfsTPxaeVHTP1pbBh3jAsMSp8hrVU5HbPqCGGa+JNHzoqsr
Vn51pwiXTy6mgN28hIIvBmB7xkgWydgadFj9F8YbcSirOEwGBu+5ofamxh3T6EfXDSjl/6lgKYqA
1mWxYa2/R4IKCwFIee1TBZO/UdWEhEGGQraxuRHNYYzBF9ZdjWw3m+SgJVqUjdZX7ZtscHt5voJm
q6iNgnBNwD8P4UoVe4RiI9BgUAvS6nxfEQYl5nrG72pOdsc+f9Rw7MnctL7NlpO8XpAgLsENn/82
rcCYnQqDHWMXQs7cJNkr0C4f+oyHI0C+BB67sP8VfPUH5/w84fLclZxriyNxYQ9A2/PhIHnOzcut
8yihSKnp9DH/DfkqcmAHKwpDoLYql9bO6TnUX/+y3Ldp+sVLkKQ/hZlBNznRLF7TruPB3MiokwJm
Is9d6xnMQJYFqbj/uzyJ7wehgVTl6kKWFkR3yUL+/LTx1MKcL/tdO8ApecB4F50Bg39j1I9e3U80
ayjw0lRz1ip5bgygwhAW/64CXMubwIiNkrnhMFTfk1q1hSnqyC8E+2c73KRcAWATzbn3izveaHUH
koZRcQqCfOY3l5PGaTV+vObzabtupXr5UJAhDFQ+6UkUVM2EQ7bEUUNvBa9ysQJ8uZa3TQjtC323
54VFuJzgAGudawxUjooN6KLatZ55rQ5JgzqX/KW6Dwxvqsq7P0fo+sjTvccdSvc+wzyha3RqWt2J
jRFFBCfgASUXmwtigH+Sxd2ttyXbVUjjO+MMxXWjXsTywPSgKcHRNszn/a69+/ZtwJ42t2JUH09f
zSPY8lUtKPc/RW4ixCL584I1i5WfJTPmyp4uwSj8Mu5N3WKZ/oAo2z+BIZKBrOs5vlYgsp8JrYxb
bLTpiMHV1u4ejNhxHgjNRKBT+Q4005W47px2V1qhUl1jG6PUD6zuS2W8N5WnHLr4jQVVkVJFFK4g
7l5U5JnLH8AkxLUD31ol6FNAKa2sZ9mCi0eThmk2PtwMhDzrpum6E7WCVVgPp775ymxTQIUpJtQC
xuh6x76GPxi2w+V+lKBTa/Ny9u7lOOuF4RHPQRNk0CkUiC5OWYAgUYMNsUHbY3TlW/uraxAWRipr
yVVek9DMxT95VKTtZ4GXMrgd3WtG5vjzj4ZN0cVKZqJO8xWch96waNKeBHY5L0ESRP86QLLvi2M0
G7Cr70dn32CBW0whmXYGbfk2QkchqH3oXXTSY7j1zthQduxEGCUdAC8zUfGdLcY8pvCZ3EWmc/X+
g/dqPI8czJQqnScwNRl0Mg6bvg9V2bXow+oOyU0s/RF34wsojWDPLoi96V6aYSv/1l7J7KMf+qSH
WwLzdNjYlv61Yaa1re5OsXjt6bZb/FSU1octsY5QpmBqxvJsFNom8nSLkFj6UvtlBddbXhZ7ayg3
z2OSt3Gyq732NCchvSWsCfuO4KFIjvsANj4v7dhACV4OJ3GZ3DnXdAfWK2mVbh6wnYAkyLzWhzzq
acnV0YT/tqlWey0GRkx0bCKaweYk7bBGqXkdWuv22mWsxAXrMhddr6QXQM6clfD/n3w0TJ+SeaK5
AWLMjEWp25DTrVX6iQE9Gqf1OJZHRSs81nF8j2Xv0WoSwpgMep5llCVwqRekFkEgZgi9M4LWMFaY
TO0szZtxnX4axHQJihv88aQDjS5eZJut7xVsOpAEKngkowtIUZBHmTRfEeQuYoum9HFRr17MQYBQ
xDZkPsl7aI2QmyaWNakPt/iHAsBG9zb74Sq7WJG25MbJAU0XtOCeTVCkWL0oUMQwBxF+0Siv1qWB
YwxDKVm2Geh756KVCB2NCc1/DkzTBfJGQjgIiZNpwWuXLxseYtIkA5xj0WiUG8US8F3gLsJmeJMP
VomKOXUHgaO9K6qUr2FO/qTw17GOolX3Jfm4GgYFWYcixnwzYzzOrlQRxxHM2wR3T86qdv0U/ojy
zA+3rL7t5i4slapkpwCagGMm7BpD+PzVb73GkYN+0XeltBBYnUSjIXz69/rE0dj3LDCmIPFb1l5r
yTgXRpPOLVMzUB7wsAbmeJ0T0XT/2vMAUoNjpew/RKZeLysRAGJX7n6OqlA8R2C5bZTB+yWRWdiO
xDVs5mJk1aGuEi/KprLSlUj8coB+CBdnXeupvDWIMA99SyQ0jOlTHljCS8DA0sYo2kvfy84jIvjw
S0V5JCNcmIQSS/jJ5XLVPqqtZvLqo+KI7UK/Xr1C62CQXm+FeV3Nw0FXrqiQFUlnV86AGgD4NLXa
US6RfP8TsIcurHbMH+qDDkzgo3pFFg3vI0aTGYRlCnL6ZtF+f7VnQ9hJj3dNJDXw+BACQbz0hO+c
cyvw42XWrKHHxxVB+SgTfHkNJTt3jI/uBFoZa/Y3E8a/LDwVzaeNnyG/1+0l0958IzZUd9nWLJLX
6ZIOZd6bJ1KdJ7FR7oejwFUuDG5NbrogNyrWt8xzhooYtnlHAMv74OoZs5NXeN/+1FXOx/dwCCIA
KpMN3Q2xUCgBCU6eGIAyPveMgnVMk+2UKrEkXSExjBpIqoSMIz5NcOuQAPR5zh+Bj0329MRl2x6H
ikGSQc2CyaWt+PPfbAoeGwy7NqZ4T8pNb6gYs4+5W7RTMwjErpwdpXIm8Hkx3HHJI6UzzeRdJXTx
kZSMy79gT9/okWAZUoLqVKjwXxP3vaHUbEKzWHqlqwQ7yyiEtiOvCJA0dIPC8G9P6Sym13Ne2i7u
v/dvH4bvOOUdplTYdZcT7q2Ku+Pm+bYL7291xXXNc70KEA2jfDbf2fqv5mdBafcHA6MCQLl/vGBf
mQ/R471YqU72A0dygn5EpkD7HyTSnbN8Y5hnJrVstlufv4J9t8pyytNanNDOOgE2inXFdXLoivim
g1CTblwDDTeU/KgjOLwSDwTKgLKOjg3vRT4EOaR/Miq56oP72VODLJ1lHN1m4+f0URxZkEMqV15M
/+eN1xg8RFqL3CWLav+bDbfJ+4fDnS1OhRb+0oFaagTw1EyTpHioIQ+ms3VDosnitwnIyKZpHnpe
PUYgTF8viqsBxEw+NRZKMXoIcwr8E5ClQ1Olawo1qmRqVUDA9XIGkkoh0M8NJZRU+nyfFWhZcZS/
Ct4DmVqzNN588ssNIXl69nnxz5vmlR+riOLVTc1oOz0/+5fGRJvPV+CcCaTFY3aJfvZjjiGFZLwz
uWpov3j3lix0Nwpmjk9/Q5rwCCTbCIJX04RS2ygbcLOUvCt1cAOE2jZ9AwxO9e+XfkCK5vC+lBzV
M7YFciTMtholyHg+uE9OBZavCgOJLCB5YxMznrxPdNTPd+DbERp72AG3G9pCI/BuDr3Se5MbDUp1
qWz+uHcuouW3lcdRM2dxrGLKMps8vMRTZERsSo0CiGM1JMCWBx8nvBrqkcJwyw3zjVQKnKc4Yz21
gU7QePTPZLxG/Z6Be8z9AQTYI9c+cZoyYNjjVayGQ6OuMOymlKmYlpsxK2yafXXI3hHRks7A7zpl
SpoycDSsFURCDOJxmL8Vcdb2o86wH8pXZ70wh5HxO4ooKx2AFt6NTu1RhjQTo9HAs6U3IX6Lowm6
uFUtHMJmHgI/wDdULQLPiSsZ7zGJBBagJ+Joj6Y9cX608pdrU3acDmhF9hwYOMolCPC/EMtau65m
aP4jxnlO93eAVLMINxJ6JWlwzzHWfuLw41SHXUQZKbMOcoIMjL4VDYnoFlTpZS2tovQdfwBJC+oC
zAMxHNA7d5ADC+RNDHdiv9MWtrWMkQMwPEUlIUiXJBBG8sWmbr7ou92sA+kzfjRuBgJotOJwVTLB
uVrYPwlEnNLoTdhxA6GOH0Il0yYyK8LDGCj3wTKFiqElPOxT9Rgi4s0jYA7eXg55LHVYgyvi/aoX
5a/RFEyzeGqmogwaCGxMPbCAkTlpTcGWcl/I3vVDcAyMhNLkNNYH7zsHhSL7nuDyf4H02cg7nUuy
d4aM5jSzqALFp/KJbL2Bi9vwYbkQ3K81i2FaWaiGlLzR7jUPUGf9n7nb3vk9ObyJBA6Ft9CGOpJl
ZdifhXUeeiPT/iVUFmBrJKMuE+mWR6s1URO/uh/DE2Wi46pz8IF2jYZ3CfadI1tGPi32mATdIETb
uagwsIdBGBYsSGKQ/YKf3TEE2thzfGbmOspw/afaNwKs31KeYeoM4onJYqyyklyquYZFoANHLSnM
hK84zKiTg3T/OidCwOmIEvGTf3873+xTrTTK0MUA9d2MrB0wgTOFVFOi4OY3zXQza4EqSlfXfMQ1
qedzPM5zag8VkjsBmOC+bCb5PsMU9QeyqxeAbSrXv+aVhiYF6vWGkTCRQ5F5z2rb8rx4eyxIP+SS
5LprBr9pAR7FjsqESD2XQxQ+PCpH2xAC8OK4uhfPI5vgiG0YDPuGC9oZzE9sZfKnIiUjEAWaqDWh
MhrDZWUEVbdApJteSYxXa3XAdou11vofHtVPP4QdfUQ+SUtH7O+Ws2z47OU0LppZMNnQWvrHXdPm
wdB37LoHszmXQdLwW0S4Ysm5C3UzXNlBuBRUkJeWEfzue6y72FEgr02uEl68dUzeBJS1cbUF/yTY
VEsibZZNABc2keoFsQdNYX0byRIqlafkUddbwdLkNItwsLGJMFvlAHwBh4h5Hdd9kuYPjWmjpo94
VeWnkSK0AtpOUHOlRvjlUWBEp3Rg6x+TjuenTmmlqcmtyE/XosI/TaOnyZNE8ECTrH/W7KMIcF0h
8ZHWOF1tOlLG6ylH71Y6D+17Nc7cMZncuHEJ8FqPnWV4b5ZsL4vXP51sh6W1wqPvwHoCUlcomoXT
xss6W6Zq0n6YH3EU0o+uZVVlr1ESVrh7GTvTtqhKHGj0TritJ1hkyjlujMrYlbpZqeC1Wrev5KH6
rrhlGaMRk4iVa/PtFRlvmaNX+7bgmV1sscxz9ctm0WRvUcZsXP5cDdKoidIeeQBGzIr94IpmCs9c
IAYwaXWyuv0uZr7JV5N3+Ng6qcTmD1bDRdB2nt45BcCvLKM5NVFiT0jmj1syTqe6CeTqoSMVrk7W
Sef0YWwNOyxP5+odSoDH/wK2YluaQB6ZDRZkBU0rAlynr6zRwHF/efhee7mcl2KBOoN1gmj5x/7P
tSKYCPZAHCaoIpA23hsNBNVyH7lHtsi9YveMCbnRYaVg3qlVJcNwzcmhiOYOLcO2xLncFshxLXLd
QeuPSB7Rp6khcQBhZXbw35wVVDyb8ORtoKV+fdpvffu3e3kt1Ja0Notqc+1JrfKYmH//cJq5yWaU
dF5CBQk/RTaJqcl+avsvcsolo6xVZ6OiQHQSNdr+Bjoad/Tq2lh6PNgMHVLkDrny+nPUs5wn0+Pu
XCXSLBA733ljd4TEObOtLQ9sJeFPl4FZKgZhO9nKNUarx/I82/PWikCH25p1ur4KLCnl0Q2u2qvg
kFiRX7K9faoznBdepEsAAYPxvDIBElUd90OBDGw9sXyy4v7rgWytk0D881ggCHZ8/5dBmNOgPzDA
JuthYi8yP3yF35+F8tjF/K38TVghXpknIRew6CagQTdVwzuyt+W0HqJWpOTk1Z51dYkyzdeVHsB0
k4msTR6l9WzqHumC47VOl/IQThXwSllvHCe6iWUs3M9l5ReTLuQfPPD9YXp2GxcFyQ6XkhYaIVcG
bonv/aR4KEusZ55SbzBuswEOXHbrD4iKBEWKPGPHYJalHUURuCkekER4kYhXDG/TknWJucc5aobb
CjF0lnQQ5n614V5lgh4aheOUaTEQfqi0hzGUlRswKWLFRGwpdNEhAiSRnxS8mpgpD/BfZxv5JzLb
U5gJ171R1n3iIY11Mt5tKmTtsTCoA+Yv1Xekg35v3yJOBlP6SwRbSndjsC7tb3QK/ta+jrds9kEA
tGbzY2nyaEglAwwyjiUgbQD1UhUiyWR7oHVyyJ/IjQZ6/PyI0RX5ZCemxqh3+oeWYjcBzsWhVqnz
poO3Bj3nDNBUfT7qqUllloFpGNnQsKRFVdT4Ep3v6fg5SySwOsV5aUtyU8hQBjB9TGSmhQZRIvrj
yUU2e/iTbzHjzm0w6inGzovhlNc48yP7gk7h5e/o+uQsIKe4oe/kcyNU1VX8C1KGqlfvw6HeChQZ
FaKQA6zzYhMT5DiaxctXQkgYx2UUh7R1qo3VeEdbqkV4Crkwvgxn+CBoMJKcHteIGvGm3Wm3KWJ7
6yxPGRGMl/RPI2ngksUgh1Xu/jKshMY7QR+yWp2yXFD97HdPGk26Ik5ahYKAv8LiqidAid21JLmA
1YfbiflAvaekvl/l6AmMQxkNNcfBe00J2nBId+mLx7TQcu/DqKlumvKy1kpqvjHF9HEnq83h/EpB
JIYeg1/GmX7ptjjm1i8nMoMM5ZnbOturMhmIqUZrO7CWlyWtAJwFIJUdZBhoaZ2xeuPRwC1D6kJn
of40Xhox9oGY0nfXHT8TsMX7BjfgCZtyPxeqm2OgBwvt6RVuHGTaXKpctWJbgW+2S6hgEASyvwwu
CxM+VW0yZNOQ0EdppekRtuDc7LVDBF/mKQlALW+wVxudvEgwSrmeB/LaaqVwxddsCzbh72CZXZa7
RbzJEHDbRUMpO6wAFDgy+WAB9U+tP6+gJJuirCXOleLJYvxS7i5gDGI/Y+zLza8pO1iu2hsvKcCw
DTp1MZsp+ORaHgat5fwukChfDx3VvMC09DOGptrqVMyhtB/vkj+JiXOgTwi5FF7fs7P73b6msb10
JFt0biZhjY1d//FGLwXerYzL3yLVEVCnt0+Wu2haPvnYRSo5Cs3OhBFYmvn9JxkfLsRLJTj+gO+F
6YgAiUSTo7VuxiRp7534wlDFaSl9g352kK6gE5eNXpbSNTyTbACrxaqEIvOmWR5G+7AZhviyIw0F
MZOg40RsZcJNMG5k9QkV1+d/z8BOK4yREA4HgAVtR5TCY/7tcDbgjlDJuRA8hAJ0yDNyWaGJ4Htl
3PpjUi1nQVEDYyDq/257J+HTtc711eVute7KolmXa9fm+2Y5qw7p0UW4vqqmOrCq/4YRQQC4gmPI
8cqYQBobXiSPbR+rfzqqtgxBT9gWEWJc+R6EFy2WJeg5JqLSKfCWb/Wxp8640ziEyYUeva3z7SGo
QvvoM5dO0BsBPBcIFE8o4HC+jBqE8iAi1yp8nQte9TmSEalJ3ctRpoGwvPNTL+m4hIisz8hREEFr
PyFy48qvU3ZeopdnHw8p9X8pz9ipVRjwzwyUWjtUeXVGy6k5d8OA8JVEC4UtVVvr5OCpiicAQSXI
obzmMYjQOBCA0sht9UaI6WYlBWWmts9KIwV6gmqx4qghy4JuXUM/4A/AI9hQyiXjQhTTMWUF2vmc
P2XzO1hAOaK5zDBi3vGnrqCNXWr9eBr3x1nAJg7Ity+TTH+1xRHB9d5wMilUi2cQLPiHURV/GBWn
w8nxLTgCHfAULJGxqmZloiTzVYzyUZGfJU7jG/6zJWTH1ElBz3okAqiO2XPyjm1SGhpOGWVvilIw
vMbUx4ZGlHKFUMG95FZy6ddU0hLl0LNcaWZBcy2mF+ZHmrx0gRxG5/0JHJQIGT6QhloeTYFWRhBC
s3OCiUayEEK3VfHtiRGOiFPUQreiD4kUZKWdn6s1oX8ad9zskNS7E5DSna1xefh6/Xh9mTMy38oO
M8r58ln/2hcsJYrOI2Ht4nQW7TP/0r10aL+aZLETbM885607MTCPyLTYhIYqCHPBgAyv6fu3IWoH
o4DS/s5uWWFr3m3IsRKgNrCXypbDqRedYkOa/lGs5cYe4nIiLhGO1pRxUUFahYNr5t7NfagHLfej
AU0rDQFzW1vSksJms5/PuKzMVS4RzBOe2f3DnNlConKNTmi4R/mu5oU6aS8BTYmS+366IUy0U5ea
3cwnGFogqh/87fvIW+fDQ6nRKoFiMUGqp5vaRkUnk9ftdmUP3B1W1P2J5ZNO0Iq6L+YSWzWwIVdJ
wuJYVi06W9H6rRpqZqrMYcmS4rp218Sl0xB2ANc7Jk5u40ovJs17jMEuMSAYML8ar0Qnpjq1gJUi
pJEwvdPBombtL4Q7jP5lptHL4o68Z/iHZ6zLSMtXUxQLYGRhayfU9Y6Zt1VoL9vN+YQ9DqH3SZUi
eFnCurqq3enpZ9JeKubLxWkFwfWjE46lLEpbiXW1Rw6U21KcfRm7ap7Dw4v0Wrm3gPK0rCdww6Oh
ke16WM3EBbrYdlOJlyGGxNC6f4W0AK48ehcyAbbEHElQvc4Wj1xgMupJTA5bli9MbPf4Abc/ETb+
qPV2NIQ4aEumIyXM6H4MzP3xwBERtCsN+eMeG81GvnxKTDIhUGmPJ7bLhQoV0dNpaeDLnpJWHAjW
EkG+1zNAdyeFqOj+p/Lt7YCy2oV8kqype4dqIwzLReJZvb9bveJlXneZynLUPCEtk3gaxcszF5N7
3DSXGTcPR7aj5ivdhxwzxVQItpU4e1h/voMpoyRK1GTE3jgc0N+4o1+gJm9hNXYl26PmOrFS3L4R
gMaQS5yQqqc8s9R2nfqHQuvTPGOBcFTu4y7HBcYKLpRinzzcoeT09JAXhRIIvUbIBbEfuaCMxb28
kw5aoFgRPR6ohCFZe0BNO3bO+hTtPFPILV/hoP0KV2gn971LP66cCQsHdLdXRMMN1t285oUwICk/
fpag+tzlmDpBS1BcHKrY3cX5IYNd0NpthNXg28tfb8BNE/d+rOETDiUjzk7Uhv/g+EWISLrr/GpM
rLJNMk1IZsQ4pKboUvod8kFoU7L0SfqUQQWWxA5s4XscUyER0F2o6rV2vEc/qsVxVJ+I2DXswbKN
3BD1booCN3nz34jUcrqP+xGjoHs5lF3nbmVxirs0wOxOv1EpOXp9xkkjpQWsb+J13IMixu+2MfwR
VAAYBBn9GEn5xlqXWjVceJ3eHiUGZ2Pgar0N+9/tKQ1yblJmz6KCL2SCRFX+ROXnzF8Ay8zFeXTj
hkfwaR1waocc+5joso48NzMGxJ32L2dr7L0Qe2J3X/08IqArwtXGvDAT1B6sOaV8r9oJ0hXvdPVO
OyqDQzZncJC587R45yzJd8rkTnHe4NRVB1K5AFKLq7MgZ+jjv7xC6nMRly4mXE5LhBF0ihKQmE+w
vZE7w6nMEy3ZK/2lGf2uEXOX+7pupJYn2FLIJaJ69QAWlxxPCcx0Hzsl7RIQR+s+NnEZjxx1SPqG
8jYDvSplxRq+gwX+3J8ndIWePv/mWix8Ryd1BnIDuOoHYd1H1YjYOzHmoDQwpqPlvpxNhZbClWsK
ZokHR12pS3U5v7NET6vB0xLWdK/PG2eAQ4bnefbUnX6CbTKJj3f2Qk8XfwnYN7BlzZhCMNwp+gdc
e6oTKHUQJ6IEaK2oXnlsf7vcOwFrw2RNYOQOgGYIny9mn4595BL/R5hrI0ho/w7fZlpE1SJ7rAFe
iLYcEfjkJIC615IVwrtzhcXV3kTgisbQp5ZSZ4fYnzQ1dOKWztv/kzBRmc4151e2qHymZpTIPoFD
zZ5SMWlYXKosQqCLakNe01LFqG8ufWhzjfBw70yphc0885zHdDJg5RKDPGfOuK06wFab6/7THmGp
nDw3oDGMa7JENokdc6eMJbL2U6JdkecoJ077Yi+VIAMlDLJ8jJ4Dy9MjQNtSNV+vNf1VWEseo/vX
evgngyVFXriz1euFEKGKgmNSpM5dbVqdu+SilgdPGbsolRXAiWgfcZhhVHP+qts3TX8tBK3Yr1Cf
zkbfAazmYembdI3ebkZPz666CX+PzUI7ZAAATQ/MO7KhVr39+cWLhozfL/RQ/q+KhPXyqAg7Pydz
dXrUuB/JpSnYiFF4FQgrCb3jou1k+Az/Yoyv8eQoH5heprQ+i5FxM/+yoxn2+zBW8Iggho5nhIkb
dzkv7TSdMoVTou6Do6XKb8UigQ9xPhvM217/Vc2dluBbzb4NWd6HY/1qXg5PJcWWFZ/uYqSN0KM1
mqst3zCwL5QbNqVTyBiTh1nj4gF/5wed2isly4P9OISP0PzWNRv/jSQCkjQKRTha7AdLKgFB0sAt
z2DZXVazMKrrGe8iBLsfjPURl9L3BKfJdSosmg08250pdKcAWCS0Aq3ALnp4gQngWTdJlTpKLkJq
h/rBZz+z+60wJu4KhXn6FFYrIix2IbY+qHKdK+FbJZmTCLje5Z9CIWWQIXqYNMbbqpZTaOChD3cR
3XZwaZ+2lnKSPhlvX8VahMjksXv8q8zzJKoXoHVJhPLDlaH2OyFdGy+WQtqMPIKstOTmqTQk50rY
cvWoelCr++Bv3fynKW1u1emyBO5dovziGkJf9M44BVqi14Ao9onQ5QRBXWahDSzTai9/JSeJNKrk
1ASTe7BVdb3pR2u38/s2X4q8tUmyObq3DH+HDN9H860y+PBQks45nCVds2MW+G1EF6JWPZlS7ROe
Pcim7YiMzLNN6tCrzPuEww7LlPybRZ0C+/R3n5KDfoku02+ufTMJRHzRfh49L89+L75ll/K30yIo
Un5tjDePPPCDHY6VzCf/kUxYNdnGxRFHOGHynowHCzz3YMb+Xnx1QIn/JlvJIQCqIP7u1zqFPfaQ
Emi729qSTzZGozLYSGetx1hjAUfjrqFilADVyatpt7xXbtdEnra3HB+/3zD3dKqzs8WPhbaOTK7m
POhbIQ4J8kfmcUWnNulzzhmRoc33ABb0XU0peHQB361UMmsyuaS3sh6ujUpf3LinAS4bOjukyZSy
+/lDdAwzhwp+2Bc0d5+PVdtdj3DzabGFery+8unPk9xua1uTTDKWdGK90KFgN8yT2TtyDggLcReN
dhcoR1Eulg5jBt978ayfp3ominNlv4JmZCUJM7k1vnuooz+rtT9ylWTtc9RCJrieSuGBPOhtAJJ9
VtN2BPkpfmmGpsz+qjY4wQH1CEQr4TtuXK4zPsEXSZrD6hEPPZoJuAMUF4VAE3blEhDzWKE7vhmN
qjC6YkTz+Bo78+uObGmpekiGEVYx7afS3ZFwDW6dhknRLmpK0RvcxY7zNtOCr8MjjyhRiYS6NUqX
r7J4kF3fjtqRExF3yqE8Ow6VwWV2wbbTURF+lH/tR9vAdbZ3+VmIqlKvmhIJNBylcOePrMayWYx8
mzE1sbMWDmRNgs4D32mm2VkFfADaUCqWmqMZiynTD64iv/Q1bRVKweiM+SFfSuKCcRYIrFvLPvDX
Sgr79mvLxxPDxicPH2CuuhjGBSjI86tEI5Y9eQqkTq5CJ/payZveFiRYEP37xxfIDsXJ84TRCh+2
5QeIkcbMqJGpx3j3SiIlExTYS67Qc0lg+WHvMqTdqec5KEnl5WuUyRrRIqK8pZEfaBdbNeb6Tw06
WUxgvnzd5Wql2fWEv9/SqUw5yWYeMSHNEz3Swv/jTxUoY+U6p4iJxrhXaCSCN1zZHSvn5eGCfS5z
uwbcrhYRT1/RYQjxJe7Mk/O4X34AtXXPR/D33dlRtldR27Fs+wFV2N1j+kGxrwpdO5lyB7FY66VK
BwaVID8TrGvOOj46xGbkCM/mu1DXph1RT48sm8zFaqL3sZZQnfdGHMT9GusbSXLQPa57kE6A+LLV
TQLZ/wY1BhCGmDhU6rczGVPW99BUfeCwfxwnr320swbTF3wpVbUG9WGXDJJhP2/8glcgs5+HAXww
gUrcAbSTWfFv+3XO4JQJEctOKsr5oQprRSY4+9SeGz2acUwuU7OX/90L6Y89kOb3at9awYjciAjP
zy9pABYwoJryqcmf+egQPDgH40IsNo5qXdzc+aEWQFLqkBOtT4H+mzMoZ8DYVaoMGQgOOrGE+AuS
r93y2Zgv8XN7GUxxwuVQCw2T3aobWYBAl9FcCYU0vbwJnvNbcPKTzDD5Yzjyxt0hBOPtxYC0B/Cd
NCrU+VGTfF8CXCnNbCa3gS3LDB7RK7ejR9ZsX7esmebuYnZkid+SZBjl+vOpjNjSQ4mFGYXs7wzz
Qbxq8lln+EAhHkgxohsbw5NWcB5PKONtAbtacjV2Yehc01WAflJdjp1CWNq8PD1uIFSDM46YpKqO
3VmMlyB6A2lJmlkiN94pwhPyuSQU9adWR0NA3Lc02wIH+XP1BtvL6lPKjUoC6Oz4OnGFuA07HMtZ
OI2/x2QAVfH6rKJgvyEutJnpp0EUaHRB4zXq/ynf65qZU5reJdpQCv/2xr1fXJv/H3M1gqkvceKM
ATjG8RkR9ZTyf+RDFML6Rm8mmSJXkKh1FN2D1xYmi3bYPHaDt3ZAdUZGNVoOreZ2Cc0tl33vXMGb
hhtg4pXYNU+0LMKUpDV/7vKocs5pUK8ONN6EBzV5Z2LTuHr40X8V1XDK6v/fw42CdTn56pRAhFrS
GI+Z/Zz9DPucK7fnQh7tCQG3xFpur10ytCE36QJhRaool+6742C6T7ZtKLBfUaX2s/JyXoj/ECuG
tjoI3nK2rS4WCViaG6BeqEK8NpKLt53CU4uPYE2PKXOrMYbqLgO5VfhmySVff5wcHflHNnN5btVj
mETHcrMA4h4FHYLQknyJVqIj3yAL0iFv4V7kQRj3Rd9Zs3qKWMdaBs7qKvDI2Wnw/L58mH+gIL7Z
waZSov4YquxIVZlGMVxBL9UXNPR+ZmNBCRRsmg3P1SuSGXwvieJzihcikATkC9tcr00hFQZWVNJR
vkU2qkODnnh6mvGAPWoJDnYAnzd+sdLl7cag5G7yZVYry+Q8gcwHwtuesw2L6saqs8uxiWHVpCCJ
qCSu6sY8paOONXKfBbEBdaRdUI8tw+vdbRRt9EYH+zJZptE8o8fV2HOmand6GUATK3Oy6dFp/fDr
RRPeHCwyX2OZsH+nawJdy8eYtvHDk4nUAVTHgVfqfKFTSXEY8/JBgPmV4xUqUyhMNHx+jElTUJVW
ybFOmNl/5DItqcM81jhoqGpFaJCa0pkYklUrNG50jCQkav+yvtRUDdjADKnUZBl2TqYPSZ6EfvCp
9s/39N4EXFMzpoX46Ll1TNBArFPU3cMmmbCM+n6LYUPXHb/ECBRdPKPDF9UfF6N+PLJv4gGcwmJd
Bz657hBwn1l7xFyXxjTaLlxE//ZkVV1b7OLFvkfvWXFtO12PSn0Jd+uZmA1sDPRu/H0EfOn7RFYM
UnOzf4RwOQiUIzBxbAQCqJOyPzDHtJ8X0O8bu+Ik38Rd49/dfAMZbZZjic6QRBAyAlZhXKLkQl8v
8SAa2dpuz24C22ZvP2apt+u26LJ1dXa5Vsq4t/GqIgEzopSVgpjbXf+lF8hQa3qNrWjKQ6JEP66q
MxszE/kwAH8IjbR9icdF/yomTxW4JYrwqCw2jgan0Cta8/5yB2qYWuUlKoosYWisuCa4piBumD8H
Z9NHiOqDQfEDLMpxSL9pXQ7NDB9zkYH9zzLWkBpOF8aqf6cQWVsA4GRHm5mCje96NQfaL9UnTWgA
0rPUsr1VETwkqzmczgHk3iywIt2pkL/4uvGKxkoVPL+TX0MMAoh6g87XF5gyKVf7jLMOwlXSMn8Z
snTM4zTRfkTxHDnGwdeZP3uyEQL5xyqk+oXlGNoHT6VclPSUCdbj9Qfge6hiiSyWs4itL2P5vVJq
dwYOePFw/m0DghZVbALFSFK//ol2Wv5MuiLcUKvL/9EktPlT3vrj6cLPpbuKijQc+KcuN5ILfPxq
8oJgjPeehL2kFuVMmnonPZOUEFPlKTXUVuTBpbhd24mDdnC3US2GLJYWLyBGcs2JZem152usPBSG
1GDXkxK3pS9B2K+yn3zyLR/7TZB1+kkJx+2ljWoTSAIFptpswJhz+LX9UlH80Od3Nz8TZ8Nl/nqM
E+e+6OmpBLVjcXbIuaHqmLTulVrns/NmauhdmSrikwj+QIWcslpijQSKilepS67uMAvE5vcwzYcr
8DdIHRBpPdS2hDnwFejKPcOgEcTrDYfo5YSkDSRwAXWEG380eiuhbSYAwERWthcSwJS56nZ7h4Fy
0oNciNSF1JY4HNkO5yWs7g+ESvjtOgddZtxiTgx8l33Cs/Ci+SeJInqn/0eOfNRA+kw1H/jZAJL7
jwGDrYizOvKip+BJx8W1/zJbsYqsL43RkWSXne9ZbBgaFFLdBSAyoj2AJ8xYrYe4N3qLrz3P9hao
ss2ezPbIG1QAI5hfcCYmrG/8eK6NJlTDfxvyMQw60KWAa9lWK5Zv4zQwnyWnc+a3KnVpP0ol9Q4h
7lbGEwLZeh/kj4WpjfYSH9oDeLbv9YxGwhzKFxHpfckaJOnlsXbo4OuX2XAKVKxY3APoN2rujQhM
XvP4uuP/2pcf/2WKScxT0y77XToKVhH+F60lXU1h1UJU6ImE3p5iws5GsWfnAS8Jl5xpKNvmoVO2
ssb1VQQuz95VM+b4LluhIydV+jkW/Y913Y1SzcrYGjzbVPNH/7ELE4VpEY6/YBDg/rcpSeSeIiPb
TjAcP3/0N8e6IxUdqW062s3eaqcn4WkULkAPqYrlRvlaBxbNX2haxYNYlLFauW29MMLiwPVsJJRc
cMz5QWMoffsw/BFeROW6rvJKOZnSgEISFi53rmeFaVJOCHsKWouNqbY9788+peEwDvHENJRpYStE
hk39kcQ/EtPFv8wMZ7+xjI0d9jFdnMXWIcqL/ilkIxtyW/VsRxlIfvWMjE9wvh+FVv8uOEy73uVu
gD75/0eFVsuRfepJfRLilk7h0ubkdYhcIqQnfh1L+LR8t1u0UUYxejb6tHjlX1tJf8Jlpd7z7dja
XHKDCNRzwk8mKq0P811QqcTNd8F648ck/tQnQv8gPIPSyNPxtCiffh9jTr0uD8+7eJYbwANa8i71
4dXa1fsySC44CVXO66+AixsoNK8QtGkboQ5idWjCoRJiz1jXtHnnomVeA3u6WKGt8SrSenHKxCm9
pwbvdgFt22x37BH0JgqRvJvghtf1RENW/sWMs/8V3PkOQpzl6Ed0rv+aHVOTNGLmXYuAUAiecboW
LCgHC3oLE7t+8bwVCwFef4EYQJl2oAEKjV2OHdABjdutA69zl+A4d0AQrAZVkO4abYXtOgTp4mGc
XL7toi1XIcOvwkPoAWShemULrtvGFmdg6S2MezvjykBIE5JFWY8qFGDx8mzHC1wHh8sY4NR5E+zr
Q+xrbFbpO0pMcnxxhTqXcIi+tHS7LyjD26QGa4s9bKrAAyuJizJqzXdVhtURzve+a2xhVDVp/heh
5CatZ66ew/hCGNjrLaf5HDceGGq2rHPQdNMhG092arZSF9Jbv+8tdB3Pf1TX90BIGd53GONKkS8F
Lt3Z0ZiMHl6RFFWVqqhBEeZ104UkcUTYea1o4GNiHC3V6MCFTeshYnwixcZVN0AmSFJg2q6TCn8l
BntA6N94axS6QU6W03ssMpzFFKB6gcTcrIfCckaeYi06hZILb+3y6vKMb1/5i5raA3miiagAArQA
LJoxtPzUzBuqdhz7Rrh/zDzl3+KoSBtYFFfFpj+s1NVHSTi9IWzt+zoDSqbca4ILTja8c4DmsKKX
bzubHABMBZ11oO7Q5xJlg+uVXx/VrKbEPIF8bH/1AeGYuZUnrLoJhdxPa1EIEWxHuL80H3Jzm3f/
/H+XLPG2t8QbLpXAJp62imALV5dm8wQHLGLU21WXshmof6CEX7vqMqWAY/6rBwbFY5zJaaNm0RKD
4tICBXuqvZu7J7KicjLVAL77DI2BcWwbRqJhI5XblZ1DMfBBXY+TXt22GM3Dn7DbZa2RIJyOtiUo
m0ZqljJlVH2CeE/azDKaPHmR2pHV6ICgvZs+fcNVL1B4sm7LgLwfCoVISntj7EJRQOlSOZsA1+vv
oB8PCt4ZW4E7SLy3crjMTPROORsktae61hfw6/WLzMKQ5cuj0mWqaCf1IEe1H72DR/xWbGbsT/8i
TEGAO6qF34ORFgtBPI6d69Jn4cOpnplUq9GxJMsiPqFgEMEUbaaqtVlCCfVcBeblecVF3iT4O97F
JLfc8RBVJawERJUabUjweZtY1alKtYSIgzcSDcUVZzv/nTxhcB/BiiYvby27C6jGVYVMpW+ninyo
lmqkkoY5Xi3D1Vs39MCQuZnvM5iRJJK/g+EfpE0YQaM4ENxTG3XBUJdwKsDpr4fAv9ERiBbA+kHb
KIJFd+JgUUZj4Lka40J5NJtWrJ39DKm7tTdRdg4rHhm+JaQ77oqXWTLtHDDmCxG0icP7VMvIgD2K
SkapbC7TmJXqxWpi1rAF1Fx4w2DLoePN8VDrYbpgXcNfH6/PGXtJfVEJ+H4230sOMpKrHzbEzFEd
0SHKxyqFspIYUZmH5uUl2Kn4XtVmE3/3ZcW+9crY36rLitL/ZEyAACJ6dj3Ve2aLZJqe1zlo8W1y
NCDEL+JP3OrJIgn/jRKn7I6ZmtAYApIunE61CMVdGky2P1Q42VCsCqZpM9ceY5qvpI6Y267N3b3k
RbR30AOIJY5HwFZPxPIJf/hsJ53Po/s8irzcdisL83niBB2JA7p/CePfKDqN001l16eaoCHp2d17
a1Ms5DPmRyfKG24HIu65xFMRY5Uc4Jx0FyulEjomS6InbZjMh5PmtILhZzF9NqrqoFaWZdCSKDLW
R6CYRK9PGPp5wcAjw/5S2kXIFirLm+8U75TFPSwFdMv+2v8v9qgBRCpjBCgwXau4SgBl1M0J5MGY
DSp62CT55j3dzEeUD+GGMiFixXBBqo1CsJXN9+oMLACC08L76YvAHMtQe4w8mSnfiAfCtqn9Fz41
pvqr651ocB8hu6HynN+ACKPYTmDkqBRGt9jLhqAiM4LUR74CQdDUtkPsbpDLBnVT4OCgLSbITQcA
B+qbhb9KIvm5wdLg/kBbMqUkzPXF56mZinWF/UPj5X+3n2ant0QR0+E5alPDXLamdoXit8cjU2Tn
eY9hn9TyM4WescVb5YSElWQ8SdR3AM21SMs0tHTVvgCeL7DA8jI18JnryHWMxBAOVj+MM/pzVyHk
JWGXRFGh3CnAw4UeoNMn2BqctLEUek58HUgjlunhSlanrcZukSOlHNa38oK+HF5AD/DRZK0nZTzr
lzlNgI+X7tnD3JC945AEOLj1IJLgBOaPvqhdDHTOGOIk57szBPW6lwKDGOK/9gDr8ZVcOyFnaWVn
iam7G3cwefzv9zhLRb2JnpzzwlR0qdISsFMWRIQDLIJoFDiOi8gn303VZizfvLw+X/tRAAMfNG3j
t5D4lOzaYzjNE47QJaUtoenHprLa7gIckls+YB4JXJEA0IbQbHARbhTQtLJq66cbITTAVfuVA12T
fIKkMmi2PS61ef069Cx/V/xwkKndimtZW0/6+axqUyxBUAkrNt1LUaABZBO/ZqAOQ7KCYZkEb4oe
pOwt9vvF/brikP1LzvkW9yJTkjQ3tskDQjk0W3MMRQt4QbIsekAjRHLurdfz8EM5IhAzGFK+0pN+
GgtFQRWxPy46dV0Y+rGIHHLTwrMB/0WZyK2dnqAoLQz9LBrL7fSM0EhvhgM7dv3BYwS6Gmld/FuQ
S3UmhpHilhoj/418wZtBzeMzNT3dK6z9cpNLpxtkJ0R6AqrnjP8sewn0UiQMnnP+6jGHYgb4eFsD
pQhoipb21xcSLMPj1+y4YS5Ii4wavR6Gy3p4a7gTN95RHSfy6CVeeEgLaD8QQfCldDLDqSccK0LH
kjNGXYNnkIWXQlNVt2py2G1M3qCuTmAler8wIPw2EVfxp5iqybWpLee+TBZwNs1Y6JOrKcNdzIHc
t+lluDf54fhNJ5qAX3rdRfqedUwAbMeOh8hXHlxBJmG0NHhmqg3JpBH5KClF4z5EqhbYajB+oYP4
g0oU0JGLksWzQhS671zLByJ+xriU3c+VLeUdxfLb2vfd5FkzKzIcPcVkK0r7bSMS+H4bY5uF9m9j
jtFgKhys8TpXDXK4vSR45P7ou54lo2wLIIjCmr9CHn+pI3jEbxg6YfIALLO5E97xX7lwUY2bRMPL
/dHidaplx4aJoyuXGVaHtAb1NGUiIX9iuNeyqlXiI2jQq7UHVl5m9F+zGKx/c/97esCqbvI0Hu/l
hs40UdF1Q7URcLAR7a/vjUscozZbtMYrOUWzNldq0O98jNTqs29BVVdBRqnSjBFaHkxr/BNseJOe
o3MHgWSTNFw459zsW5GOwMki/YMUJ6KWYQ4qR2urZq+vDsTOasD0u1IHCdQh4K4CwbEkBPDzq0eK
pIuT0n3AZ1WrgU01cNuI+waZ+dBss5W0lWBzb3VOejK2owrnAKHg1YfzOMeNOmXIMXl9jy9P7i9v
aS0RpmICi8mu+EE6pQGTkIMTD0FAkqTtTjtoqP+kvspF9PFsf5AqL1AOKX2JP4CXu+NbdAPcMtGg
w15t9pwuOuQCEfLFi+cQgBv1aZrLidi8ma9w6eFL3WPEh6esxSDHqjm4sZksynpIGrAgSD/HDW70
LMS8A0zYt97IaFdRmZoIyrEqmlYD/Xw1hVu05NNX9QbGnlI0LtxOoDC99E9FOF0QP94blAJvK/+l
pcA5iUu7DtiWWQKCNERL1HcPVmrPQKpzczrSiqRytC8GHlogrkJA1da6ctQYGc1H9sJ+eXz5WfQd
YHrjPfojjgOAYH6h8rtG5q17rILNoybq+y5Ehdb8w+tLCZtE5wf/OUOy7HFWdjVxZAk4uBfvLDy5
9BKT0TVV59R6kEUi1RgWuAOJTK+I2ispHcVC06/9t1iypvvHOoCI08bRjYAqUtGGNgX53eXZL7HL
qdvI0YGjtOJ2kasNnE0PR1kYtyq8TyZ0eo+oxDY5ordesIiZS11VOTZUmYl/Xzt63lX81s+ajk77
DgdBWwue0DmyEAu9nVpN4G2hAO4tYTYByCDwq1k4HL3qYPn8odfJFLetjFElilJm58v7kXCrgcnj
CqfYYqdgkGzM2P4l4zDvaBI6RaV+RnLyzMLfUw1MzuV0hSwE968crjJDj3c97tQ8JnUYj3fX8mL/
s9e28CR+W0YIXLPTTVfl0UuXESQ4eTmt8F1LhxUMJq+SqlSn1eoNjx6KPkOMDfoePhf55MlewQS+
9J2A878Z/hycYRK2unFhkU/NVg97oidojF6+rQWMv/qYApkYJpkZpJkvgdau1Mz8suuAaisJkqYX
P839C3nw57rXwlGuxodjFR8ac5+OEhPgwNFsYfMJhAu5IqqA98rM4FkI19TBfGCWl5MwqlMtXnRI
34IW6Ul/riwPt052F3dlE0XKq7eIy3b2d2Qk+h9209uAzvMjsU+vME9PBWp06ZSKJ046HGc8Ftmh
f08hr07/UAUfa5SGnh0zQT+T/icjsrY9hihu7cvpmd8AZL3DRuJKoMY4AB7k9lZm+IKuvPVKOrYJ
c/8uba+ZUtKZaIzJTLHu9VyyxSyhhJF5nigpLFRbbHBP0NXpwZd5GBIlPoOVGI3sQegmnRDC+Mja
bmbcpZ/TopPU/Pu8KLn2A+wUb25LTPzIxkcXn7gJhLf0382VsT4hPx+BL3ZDE4DKBet/P04Z1sJQ
zSXmu6Da0yPsWBESaBNqeKmUexYXsM4b+1zaSLGO/Hy+VvbfnzPS6Vm+CdPWUbD3WguivKATOpRg
wfuEoTzKVXUsAhD0yfBqp+PsQv2S/R6McLupOogVH6vFEE9l1t3ycAqo01gPVW1yTOfIhu7xHkl4
pzu0M+dO87LUscthxZq1ZuxjXvUT2QJjFDvh/m3Wnvn5kM2sYAwzatXe/mJQKa8jTZXYFokgVxsW
vD0CzUD+j8sUX4q9gYHI24nTfs7WAnhqiz2vmC6SY4/0vvbI2W4FzSPUwL0UJBhi2fEPU2MAaspv
IZZqAkdO/+MS6VxGd7HJwz94TQaGnMRr71lUzo5bFo+SaaRlzOhrypTRfTJRX1hOtlTdR3m+0uPs
dFXH2X8xat2VIG5N5GcvGSESVvfvIfpIIp39Fm/JOL2eXRq4nenOfudnjvH+0wCW12gKLfWKDpID
iK3Q8DUnjnkr55e02XihXFHk9vm3x0BstYW7JuRd71KZZClVKQOEASQdco6JMJGRcoE7j7FNWQHY
yDw2/EzBfSc4+QouF+sK9ehk68jVU7fj6IerzAL0rynCitM7XiUltBxLAFCZVpPNl5YenD+eZPBl
IA/lpyxCLO7WZdgu4uNR2nnOBV+ruf5SGxRABSSxJ8k+4P9Da1Cg5AHX+fpKNsC2LTnH0jJpElhu
QKCM/ygaVi72zv3+m8RiusS7fCTA03BicfnwCAb60X1stE3kEqLylpti0IpcumtpvozKJwxT10ao
ua83aYAAzPb8z25jhpDcXYXuPHWxT+ddhrMg3JtJqcBb93vARPIWkvkoDd9kLnclqc4Kr/B0D5+U
4wBmraIZHrnF/UeDhR8l52GHY36oLlok8PC735WOaFQRzsxwYWsLz+Y487WhvIui8hN/PPynmsBP
tlQ3Z2CZsTbNXnDOE+HIX7NnauA0nSmiEZycTTaZF2wF200HGNBeJqscqpyOzS+pbVUfvF04J+N9
zmEgRQemuwgEET9eQU91vXa0DuCN9dry3mZOetGttTRlIsUv0pm7p7mO6gSgAraXHix6yuYj1+JT
el2xAtp2jpAAW3eOx7TUIIh1EhzYqhZKqvWRoZRTdAbJjupY+012IoOm+/Sb10/JWbOZ4EMmXZG2
hhpsBO2SBuWOUQJHU4QpPVSmDTYhKJIZh/Ar7sXm5SQm5r2L+Xj9AllJwua6gsGneQqf9rNxsntx
6HljgUCkgi0CJN3RGywVVN7E3RuIFxRwaOlUNeS2isPIgbeTmQd270LfrodvFs36WMV2xvVyKhwZ
v+GKNN3M5K4fN1ta72xBZ+6gjQHoAqcreYmcvvsEUOESQghFmPyRogPAot8oxsXZBIsMUY/Y2vK/
NbzbLt/sCihGu9IUXUbEfc54s65ueGa8AKy3pYWaOHB8lA7Q9I6BBQe2UdGnfN+cEbDte2ehFRHy
O6tgDSL1ytcTgK/Um6P+LJgZvdgtG6282r1kSEx9WyJIhRTX3z7vhkjmgk8lBqIvPFsF2fVOQyFM
pKabZ1ilbtSeldTS2U7ZDY6rvgCu7Jf+zQ7ytlxtrRjJt37e3QSprnEGs3dz78u0D3eoMQj8gAeo
Fi/nq5mM4ptgXnDOaZSeS2vUTosqWyFKg5X4DQTcP8+cLU8OFF2PM4nbP+ALOMcVjxVAXLDSSXAg
3wLwCxys450dimK0R2Zl+nuOObIhMc4c3rp9Fw6l1bWwis/7yud5kDgCs77bml2Dgwsf9O55uhsl
+rqPNFlSBTj7tkb55QX0kkZRqRL5iwdsTLWViBM9Kv0Q+R4PeP3sXoU/oWfGyworXXGPGyZ2V5uI
9qAobez1GdwB6UFGO8t2z5vG0g6u22IP5sn+FbA1SejiHD7Ej56sPe96okmDV9FV9n3s0CZ2P5JB
WsdZJRLDWb//GH44fHx62hU9n8BhX/Qf3VpHDoKfy5BfOUds3wOpAL2tbtwqdew0aV7jaolsXnmM
sZhGXqtVCqSCzXqat9nTQD0ZHYy0Qpng4YLRvUjjVJlBftLGupl5Pjpx/b1HO2BzebAz0aWmxhHG
Byo4YqI4vKYGUKJzaL4wMnoFWpMFc8kM+l76dm1MjADELXygx250OHq9tKt+q8dM4NX3g+WQyLun
UUzSlqXOpic07f1GOtBs/txnPw78ee45jv23a2c9clk4upZQ61QWhRn6rCFA7pIEYDQhk9gzHjzP
H3v730zlFG+GP19UTwZysROt2EiRfEBfilTVi+4cfoZDXxIBqfhyT8xvonwFdFEEHK4p3sR0PRAy
3o37W62OFWXhFhU/Eulb5aC5JSIgZlt8e9cKAlrdOkvEnwtwOmL/ohN2jGHhCKC29uxzNmPuZd15
1NLAIKpsum7Xw2QNagz7zcf5idIZbZQSpNmPi0g2UMkucphdEOJfIxFzm3Lqatb1hOmqeySzSXPv
Ayt5Mnp3xc1s5os5BR5xa6N91c7qtBre6/FZe4OPXv7ZDewFXWQi3U8v+zR50LZb6nf3k6i+feZH
1O0ET+OhZ/j477NBI/yB/AabymX1ahDj19JzDNVF6zgk07eAmjPgiKZEC8LTrTMDBeHp1FXn8pg1
KD94dRNXGXG11OaRgmd9n7tn95XwbEMb4/azuDzMc4m3FzzW28WidLmNrPFE+mda/LpZ6jF1xCWn
SoZ1kYQyUw+v0+BsD1KMyVLsRLeiIBxbkojt17stW21QrkOcDPde6L1Ve7SZitocwlGE+7fdttJc
SUD+LIgHvd7e8EWl17AIIX2odRMnTMEmTQQDGw5yOXx7jw8CHR4oXqxKkm8bkz8YjSUU+aeNtqxc
tg/BuWzeBJJyhhkLkVo/iq5ZbRVjOgWDAjrcErkvtHqR9UgaXzt20YSg4ub5Eh1IY8Ui2WHUPtQE
GYARLPVOfeLglVCjk/4rs1Q1gD1zam7b2aGBBdv/EV7pj2DalQONTJ/bbCp33ORSFqqasakqr4re
uHSk8y7DNkcmAwaLYF7KpkLvah9fwMUyFgdB6WgsJWBkNdiRmUfdksS4DkMe1mg3IdpIkqlhldf9
rK4hZQBZSrkQZDB0ajP1yzDBiml804XlQdx2SHgjRkN69JwIhmii8/Pt1eUZwUB3dQE2Pon01ULB
wobAo1IL1ie+KOz+4NNhgmfJ19zk6n/2/wJ2E65tzt3zw87Z1NVRzJH0T/9lXJrZz5zfTqUD8GUf
f0OoAbpw3BLtbMyJfNV/7br7mkCNX4E6dwlUWM6J6GcFV2HXtRaQlYVij3Rt/sLVPskBVAdpPKgH
JHAnvGAULudrW5Az1gDjMF/5cHO/8JwVaGOsQ8eKKp5vkTiXEtjSxcfcxQcWp95G5D9uLpK2bs/I
igIWjlO4DrCnkIMU2FCoAh5/wM0UEPY/XbBj9qHPDFTwjyeKcBZZCZS9GMc4Sc933hCP8JoHvh7h
KCpfFtb7ZXW1huKVflbe+9UBAIHMYIx58Q0XXf4742KMIwNc4UBMG/bVvnO4ZRC4Ww4Leb11oPOr
U+J1nnhoaDzN4yb5EXFTq9WCnEAQU8JQFd6LofmEe3kVWLP4qc1tJnxSM9z0EgkjxPh0Y9jXIXf0
ze1RLEkvZRC6KdQHsXCULzz4oeovs9t44iGYDCRjEBlS6uPNws3CVZjo/5OxMX6bDrn01wrTIXq9
t6YLysajReh0Ns/SctzPy7G5MXD6SmI3nhnvxIrJPBlN1d25mEUk/d/RRxnJEME7xorT3Qh1Jonx
YWFbuHaq1abCFbsOv/JYNrOH1Xk4LUcm4BROu9LQkTLZN/drur1hwD/t9TO0ORbg8GthQLN51Hov
HQiMmprAD2n95p+2uWxpu+S7JXLG8mEtCu8rYbETevFZPNHup7rxzNl341BPpsHGqxBDTRRubY3y
0OW+ircLlY7uBpXltt6g8jkKyUR900t2G7XD3/pRx9l9+u6qEvRPNgtPHWcRVM+KM+k8QNHJakZA
oBjcK530F8hmNI03v0Vt0kOc1PJsFwTfA/R8q32vy93bmfb2XsZpvN/HRRv3KzCpu9mn3HtbumTZ
Hk1B9u2nYcLp8J57UClvu9ukvKj+ivhxs2spsZs95vJ08clpk4YFBuPhq9bP3Fp6ggaNEYjzeGdH
XIFPYXdQca8SyP/cE5FevhFICm+1NFlxPeYvbm0hvNkZ0dw80FXQdroMkMt2Cmejf00Oc1Hyrsap
sW0crdMpFjTKEsAvRH42LtiklXpYVAC53ckwC4M7LrqvnwT50RXVcOPIw56igL68YnC2zIZtfQI/
wT4DIDgxao29fyELiUFYWTbTHSiqnl8lIhJFM9EwyEXzsYA6EcLjkwp8Fi219STzimbayy94A7fn
ze1R4/3Fc2h7RH3seQyspDZTI4CyseQkdosJdkEVPQX2zVus7SmJnOyNs7Hv8x3WHzSebT2r7e8j
gADksrFr29FOIBuVrgtRaiYdFLdJXScw5bB40tE91056DJJF/Dh7OLYm2XAnIqdFq+YTGq72MWq+
oLVFipK/fi7eDGidHey0HOOdsl2DyjTBNhKFA3zApzCxyBEvKYhANZdx5033Hg86gSUCjzn+/72+
no+G7p7Y4wHuUTYtdh1tda+ZvAsn5NPdA1QMcdktitXGVtCAM02QHkogfQBUR7lfSrWzZfyxTwu6
fF7seRHl89ge1dxsmfEHS+ByfXr2LE/1Ch54GM1ZhSqvp8aPEts8YFyVwyxHL+uznMBYKdEySIUW
f/aKCSqVdJDI27lYerTfdI5KWw3lNaU+Ya1a2ALY5TspBqnmButVX5D8ZYZxxkdYs8uvKJoeDcpS
t6yPL+z0nDax6BlxomUcQ5AQi2825fsZpIWqevMmIil5B+mGxICcsMuYb2B4rpMo6DGi8VCmz1cp
U6tPIlHwxO8qlQCyJJn3vEpjH/19f9P8rjXbd/1Y3VEhNeIUV/s+ArrQhE9Cxt/MAX53Y1pNlCSi
XE4+MfFd8DPv1UwVS3Dgnzm61nBeRYmiyNfro6fDKFuP5k4t8xQwaS1JoP1y9RwrE1Y06xswIZ50
ppcwbpXce3dXvdJXTKrp+J44zhEVY9LdGQrZTzZMcG3satlumFzuaEw0B+mIeQdLlcsLE8136kCE
qJXC3E3YKyPgV3lu38T8KtCeDe5INAtDj0u+xMA6ehg3lppLwM8smN6cQTxsqwZ6PLX8XbT+oBen
ErykYINdbANzNYNMD0HbmFz0K0U6tAXM+rewlPbnORwqbIiaTTCv7X1AIeoZN831EAZnVCcDKpag
wUuZIylWyM9lgVgReIYxbhFkpCAGk3kLG2lAByWzvystCrwb5S0T0PFiXb9d1+rL+jI6YlH38Me+
V6Te3DBgskqbaW6fPGX2GryUQ4hx+m9K6XycaN5h3OXYwxdwTewxj9Tu/P1ZNCKre6uznKlImX7J
TQjdXI4Z7r9xSElXUMAJ5QfUw7jKcE5IZu+kO8iV7OEjzZfHFey9VBy0zuH3T0QmhYx893HcVyC4
ZFgUmyDCbQCUmUBhmBaOt/7r2QdkeaN3naHLyEP7yW/sL+gq9sTIrbAR3TWDkH+a9a2tmT8YSTSe
fdDJuBMzPHKcLV8W+iswirc2ar9sqMjKpUd/O+R+UBP9RC8CW685S8hrF9WYlfJi9v8Vw6QNPZVH
1ov0IgMDSOE0PHO10Li2q/t1X2wXXROalwLqFrSeHYrgvE7XQHHwKDCCpX09wjALXQZInU6hcmFI
HYTxpRmeCP+fzR4OZ/89HKdbWcwd24PqLWE3AAZt0gHzMKnXFDcdrYZiarpoyjvQUcGt5XIe04oE
YSq4lvoJ4OW18jA6SJNMO2Nc0F86XrH46kx2j1+fueGsfmKhagAg0T1wDghV6lfic9IB9s4QkYcV
ilxH6pB16M+qz5UO3ciQoplwRAZdJXTjtsCLSfIP3WDU0foT3DqyRY7Rg1FTpy0eRXyGZOlf9DWc
1ogo/X1N7TWXWaH1TrkVbECdcNAJe9pjosUVdYJRM6cVDJ4i/U4kaQGwZaMIr0Z/ent26fO2WvmN
yKPn0ULFYl/9XGlgOTRyWH40XDdVsFVQr+/bORr89YH1cPmt+Aj693/iziXz+h7td9vEok7SWbqF
A6azdB1kraXPVY35xYca1yGgCot1TlmFQT+lBDT7pAZRlAyq/0695DRo0apusah2zuq3oXOKp2gp
fZPKbFegxGG0yslS9hyaUpyqmihyaukI68LQY78m1SVfv1H5RvzcWqyIJYDbTXu/xYkK8SdmgaQF
SdtR29FPYf42F/0a8IUalWudq5c04rV/0UipOGWKVAAjx45cuupxABa0rTYqYeDYL5tp0GJQOTxH
p8Gd/Uxf7kFefO3ATa+LkLpFx/hsrcT2gKwqapdF/NXDfsZCLWmoN3VKbk0c/fNqMbymjeJMbxxi
JSETeTANFOsf50xPrYagotx0GjzwOEChwDkUK65sQL/mUQNnVvU1rwZEEGJ0dS5Gkx8dlyYC77ZS
vk1HXLUJUHH65OfARgHLdCGo5E5kTtijXOpp5a+ken7uW2klA3KcHnIJy9W5fbDf3xqBprEtImVV
UoxZ4f9zDA9dEjvJX7qxdcus+zCfDz6k16IOND3mY7y2qYbXHavIRfPMghrkrqO5Z4chCkIGwo/6
9TwFelQpc8zqxEFEB+JZdNT9hK8UCz3QMQFBENsxg+ugREr2jCwybhloU7w01LGfliYRPD41lpnU
sX5MhCXZWBfRK+Dc8OvVT0GewAI2itMDzhiFCrxpYoelebSiHU6Cn25b8R04slVogxoGglY+9y34
AsAuNJ0pb47+ChiyajIoA4cQkZrA4WfdGWZDBhOx0HQEqEOxT1RsdMJNqmWbtFCZ8dUMn2szgdck
tKkIf04z7Y1dkif0ZQ4yKwzi7D0YxuU04/VXJLboVHizsFCOnRe87g4KwiS6fgbEpjirbvA4PQt8
RCAnkREHuN6HEc8DwuoS5LYXHK4Xbo1Jrl3ozIKAXbAnN9cZoe1VWZ3qin48sS9Uv2wFBarSJBQA
bB98LFMMrESAu662ae4xYwgNi3i+cuvmXK4k/f1Q2r4jZjbIqoQSCLzRahvEKAAE3WMqu6bO9q09
4Z62e2qmpsbzm2WsNJRIxLhpxd/cQHim3JsIt3m15F25WRAPsfsPtPoxU+N2FUhCKXZfxORHop3p
qgmF1RvvAT5BbmuWTCidzmFaEVHcRyDpEL37eSrcWkyw+5aPPrtXJUAqCcNUjD7iZxeLv3QSBi3A
DV9gZHdBAn/hq7UHfBfQs2uwvwIU7wRCitptB+DROSh+Ab3A5gXO1v34oktZPPNVp7dy3g+5CzQU
H5OT1VbwFa2B/ZaQtl6TTKeUqQ6LprFcLNpdDmoZMvuHJJ8BRmzXXsWuSW9A5DWm+xZX88mcq1Ec
oFe+z5vW00cpbE+RhUbMr3eEHGeRF5UK1I/5XafB1QgwUicjZFOFywUslJgBks40l7BLu+SFdxBA
RBD/X9GH/m8R4qIcncVdFwJSCXY7XTom9g1PCdlwzaPTTxO8N9+OclcfZPGkV+7ZeacKePzqKP1I
16bZxhuUch5Pjz/a7W8XzlItzc/lG8uJcmTH3fMjuK6HM7aCF2Q0BXNFkEhXBUNXZT6RAoK/dhVS
rLLv8qcKIw9Qb8pd/jkvKrXjzOjKzam7QUEJiRCap4v1J6gDtoTzB+syS3AuX/LWGdeIu/VK7VLk
S7NYRI7YDr+yzdCN06rGpdfMYo/Cwbj873eYjMqsPFgPaQkA4hmZSq7qqwnjNUgr/qioWoayaHhA
H1w3EnKpqV+LkViaWViwDkOy2RU1ieFprJcs7JNzy7APrAW6rOLaQpW8qULpCnZb/MOg7R3JoixS
I0m2tuiDGoe0R6YZqGRBW8XV5BWE92FbGX0W4iS4/OFNlK+lPTJC0dYykcyGAUbFGCl1Q6ErN7NV
p8i3Jfe1qTWJIGdKd4emxLXzIJWsC5pHfgpK2cLTSEKLxamA4h0G0ovAF3Tf+vV/92B82Sci9A1Q
V5bDI5Ajpll2x7gRff06C9AHxKSNIPOqJJtevwED3+toogUr9OHEes4a7xMEwbGVN1NUOR8J020m
5jJTOwp/EWQg+2qwXLiIeOGPaM7oDHQ2Q8DZ1Nb/2hIkhavsxfUTjMDGFfkPkazFnbAKp2QWuMsF
NlOGFzWvjQ+naiVSMSXpZuhROBce8G9S2D09uuiaJqSkSiCZet5tG0cAjl/Zc8mJg9gtJXdcCW1l
mzl84syekguXgCFomkKdyRen/nXXXLNkfsAk9C0rpxpOkTWJ5SQ99vN6uxKSK5jcvWnJWMrhnxvK
PZWrJslbzitM0Ypt748CHroCJWreGJPY0qoU87pOBTLrbmt2j/IK8PRPuFOysp+orBy2PxCe8jRc
1keYmPe3kbCcYWO6ezwv0QA84xbeqgYUHrHfHLU4C/dIVJjj0vDJ05hgFjERcA9uRgp/M7BoqNWa
w9+NyRMl6hzf31ENky/8z/RCL27DvJKXzhWjHih7y5u+ZwRVpzBoL9uHBRJSICs1grAu1vd1J3sb
/LH6A5Mwsz6ePI5/vK3nft2/ysk7Dy/aKcpFAuUBCuNd6YJMyZ714r75+99Qazv5olcXDONTGk1S
ZAENZsBrS8nekjx/PXROO6cQa8DtfPnZ2Ev7dgmKsCkHl+p6I6OhNKQnpfs6DtwcEL7hYLnzqA7z
MW87k0JJQZ+Mf2yuJFO8AuN/GRHtfTgDYuyNSjdkfrvXySFD52HiUhJEpk1qGOewjcDMFrSS8kom
2jnA8b2tiKO66KDATsJ2aHXZmxy5yMZ9MO1Ds7RWa40CEwcWl8JXk4zSaVpE8N6w1cxpz3TECAEo
3wDLXSKbR1nQkgsRU29mEZuyWQiYczPSM5EO+Bwk8rGrwrtKLdcJa+IUrAQr+RXxjQrYxRmMKEeP
Cg8qgJ9i/PqvuUvYTaRSCKHB5EfYTiOo2GmO4nLDgX9Hm5gBbIg1mKqMeZHc5ouxJTMI7HYuuvT+
TzIbvwekL+XsGYIbc8GiXUfYilObNPwkE4K5REiw2HFwlTuSx1vCGA2gIUghmZT36vGoXrYNOczV
rWTfSpGiIdfekQ4W1Ls5TDoIqUvB4ECi+de3HVxIJ79tFnB/auJ5Q5Meyvsfzgvi3RiSyL313Y9a
CnLYPlUB6aENZWjf76SCW74/fLrqtHRaqusQ9tCL0GGz0TD85Y0vQbQdTewWqhmpTqw+NoqrneI3
4zkkgFbN3Xmc2vgOL5y0c2mwMhxQxatzrWeRGXoPWSXOdQP2euvHy7KvnYwPz84IuOKKGuchq+LL
WRwa5SIWF5XHMy11S6JInF9Vir6NA8WukCfi8B00vNGpTOMSmNHFT+w4nf+VLY9lutgk/4Ro9R6z
8CwoHCYfA9QE0BdYOX2APmneMq0V3smWpSU08IQxm7ew3S4n9QHcSb2Zam1s31d9k55Z0Z6ECJ7C
q8DUZhyxXpj4sYpDb37L+KdgVkBrzbPIQWsK502lpOS5x+meGVc3Tkkr0i9+3A8j3jg7AX1KuYjr
/yW0Xcgsny2uNK4rYPtX0XxkG98E0I10BOq5SACiy0PMr8Y35OMRW6tCqsUW6dRNV1+UOA0Ttuh/
/LOQ34UxlZKh7eZYl49I6e/3Rj2/C75p1+DhlojZ1J9xRbMTEk/BF4rxoYTyoeyHwM8riR2+GOGQ
f79yH9jnvzJpyrYn0n530Ovr2z8NSbwPy/IPimIWGpn6ll0Vr3affWKZtvSI5vsIj+4fdjDPoI1/
4CJK9HjODah8xuA1vKGoZ/bqtCCt7oSOtL1ruZN1zQKfk6V4NMFHToetul2by/2RldoCE995dT3W
3ri06MCrprkX+XJsElGlRqiERnBx0gdy7j3WWGTgVxiFi/AoiljtvnCx8eG/SWO8GNJT5DdtX2qS
2VrDz7kT+R7nFWpQN4onkz14WDmRoFrfAOMxjgQ8qy3XcaDC/61xbNvvR1a88x+fTHILCNrHaJxo
CHADxFlN+MJLxgStEimkCjIujiF7uaDyJS3wquSEEirY3ls94xHKzMLzqbyULoBBsHfHYvFKDJmu
2rlKLr3+BciNwNn9boj/s42brTc3soFKHDqm3D+xR76sWWAZ/5ePB6OX0DnDRS+29T5LMAHYbeRj
lVJT8Kr5ey8bXQ5cwunzfAqixvykk+qbyeCaWqEyx8XmKJNPVOLqXl8QP1tSi8J7l249Wg7U7dak
PWvSWlPC2dY3WKn43qdcoPdHL8rypJSPFO/Z6H0AapcNuL2yK90C5fGdq75FHwfk2Gob0mK6SMuM
odsSQObxErM9DN3H1h03QRpq5oSecU2Ott9BzhlkG0C9bvJiPaF0bfDE0j6Ddz8VvSitgztN2Arj
hTmpNcB1A5jfjyj7Ja+JNirZQmQCefJjYRd+fc+8Kgp3h/J1twD30zageO8L37b+qj412TXnF/iG
KM7hHZN4jZBXGYQ9TAFht0zmtC7pDyDbZ0OssqylWaHpAFAyxWmeWy/YC9vpOKi0FD/N7Zyd4OBi
ti0wn992NPLphXjfdNqLNMz0Yp5aqlwJNJ3QxaAHRlf1Mzbbd2i/hlA1oV5fEiwonHQNBOTyB5aV
+i93NnrkdlBxaN8tAiJn5MhuxS7FQSv+o9p4GWvMJfxy+qQnqrQkfc+aE1LN+nWxOdWasiY6yNXl
jf3rKEEnA9d9lB0/G20tYs5ompjYg4bt9hr5ujqmYxlxblO0GoeHUWZ3WWBsIRmhZ6Ki4Z5QEy/J
xJfQYGRUzpkF+6ok7SNRPoWXXLhddhPmylc6T1vGjHVa3yjCAzwy3DpsRwk8DUreiqVNpFfVG7/g
vxe50Smkk8EmEKDdafhzAXYJDuIQl3qek6i4eaZNvXeLuDU0IxzgDv0k+BlWpgtYhc8hi9MaznRx
n9CIvzCKTcL0Na5Lmsq/kd19dmKs2Tg+FUlcnoblVB4Cxljo5R2WRy1bGAS2oaXxx+MOwCrsTnH9
LWFdDkgoEA//UgxcE8g46FENFNxeW4hpYQTxu2FWOl5QCDMj1r2th3vWBKE5DWnKjyqiVsGv190g
mVGcGMJL0q0WsZQvivj57tJDvZTLr1tawucgMVGVLTjTv8hLFX6Y0j6uLMXOetLIluHnwZwjhz5I
nDCVJqCCg5jqr/R6cfJ5J06jHen3jgXVX1foyxESYvnHAC/DT9p0OcwxJPd1TSya4WJfqSljMKNb
l7choxHUkjdNfsSNgjZnIbzHGQVw8XDszuM+aRVaq1JFhK2KXaHhFZ6jk7olPj7O5putCfN5WdhK
uzGVS3ZJdDy37hZT8ktlA/NBfrARPtqA+vxlHeuhSQ2o6KY9ba92CeESAeJ5xALhElnP9YUWLJB6
VE1im8QmmfnZprE/ekaIqbNjjxtcf0z5vlCC3G6w5uiwTfh7l+gW8EJQvN2CHR6LroRJE73yy93f
oRmz/jExmS407R+epE+9GOOHQrVVAiyZ3AKIRjoumoKQb+vFb1u+sftMA6l3rJslwPo1N428mCcZ
gGEc2khqf70e+xpXRQ9FSAS8gxox0T1zjRcOMwmVZCCnVjJ9uGluxYXKQpzNtEtn/05xkAMxcFAj
uI7Tz3XJCqEfTis+9wpnFzCo0hh6lJJkwlXFQUt0Pb0J/G1Hy1UNn3qz5++7clqvioKvdjdv7aES
EJGZv+fk2D6P2OAw9aYB86BDEeOcdtdCKvMOVlfEnQxYzSTiSy7DvVdmvGff6c56s84wv0GkM3W+
y3Lh8qvJN2veRhHdBv/WFstHS+A5uMO+HXXEW23XHvPrDs5yH6btvRiyJD0CkJacx+l+vAq2auiV
Xhjx6qBVaHkHNDT5F/YfxR0Pxlc4JQcgpzD3MRE0KtxJc8hZb9Sho06rtWT6Ec6HIBFp59VlMkUB
y1smIUa6WLQMocireYiB80dzd4LMapnC9Uw10UFN2FuNv7akbw3dWN/zPkQOvCKAEoGWMyPzLv8C
mQeQxoHX88a4i3YVpA4IvSjAF5zs/3i6deKlPw4vd0M4WFXrRJg5Otf5flt6W15iozwDwoRcTlV/
sg35RJTQe9f1SGqelly7wbRJKzUekhv47zhAKL1lIjPr1B/vZMKVmT2d/GEXavU6/EZ74/5WOLSY
ajIDyc0qp2DeVSliuJehHsBNZTaNK9cx1rnKuBTDHYK3GQlgo6fVxaMI/Ue1GKBBhHnpK/gcOfJN
AUqAFKtRL4ltcNPHBrNpUYv1nVYW+U4QOJO6pw9/KqFwG7Dm2BGvsFo1J7rY/htChRRzj/O5DhgI
GhAPiujgalShXF7U0Fuqf7lZgqissPGONwL5hShyPv/xTidJC2YSmlDiHVjKj/T9E/rCbXH/3B7o
AD8T3cCnRBl8Yg1i3hSvHN3V70vJ+V0acBp49AvYPWZIqCckKHFyUPOLi4BLnkNHImCNFPk+agAR
/N1RVkjkGTvvIAukZByuogpkkwu2EQXWOvRsl9uykza51Pkh5jOdXz7kec5w84/oEyy/+6gDLRwV
OMVaeu73W/8oCynNcGX+OJC00J9xiJAopEb21umHuqui3zto/Zi9giGN740pdijMgmCQeSr0YaN0
4BF35cwnC4FDv7qANHXUYDZkBgwc6YntmlhP+bQTYdQzGl9uqbCPrTQA38c9H37W0ZFYdUr00PCg
kgfe6ek/jEoxAMo9nh/RfdR1yMFfepoqjuX40YBjmvS8wN9tttT5Q7hjqdCis2Snvnf1Iug9rqcG
IlTn3rkT83jnZ61ZNx7imsa8uGRuJAXssWP7C/96jYdXsaxdCmxc7yMt85iG30WV4PU+ByQg/SOV
0Jd9dG4UbTQhzN3HkZ4LAH8m2GjtFajVjwJxfNjN0//ok12jdd/h7QMOz/X7Qjoc/suJnnhnWx0I
8v/+sd3+zuUlQ22ggDh7rPjhK9+9o46hHnLuJOuOLtNOCTPlF4rOOgKjewR1ZXIBJBzJk0krfeso
5i12u1YR2wZImqtwCKnY5PBEask8R1gven/EjdeQsQ+UzA+/4d5qeDmv7XvA3r9qaFgj/dileX+j
D2PPTIJvxH0mt4t1PR7EPNO3Xzrp1eFa/KBIGRHNVOoUaldwaU8KyrN5JasYKIQrl/MVD/LBJJcy
8dEwKi/8ak10xlPE+z3ei0A2D5KP6Ecm900StT7zaVvzGp4QU4c6EQhLeprqo4uJsPF73wEaLljx
86EZVKWAFg14ARvdBZlArcVMGDzl1XfYA/MnYmQvfIAwYABWzNEgu9imjisVBrlZj7Pd+wXoypsC
Z4sXMTRG9aLUWRUMbm/0Xuk4FbM/aeaVWjCZAGq3hB/YvvBgQbrX9SjcTFqwZW36ENAz1tskAspX
QGXTYywKaYuGUmnj17KeXrOnKG/PtFOw1TRIKKkjx+LbYvhmttGTDIvvgONOjats+z/R3jx+FrOv
lx3GVS7tiK+HBd31uKbEgqzLALG3KmVTxswkle+U1aTOrBQkwOP0rwbfkOgPgTYAOHLW7O3NASJR
zhlYgQFGgMq5XCYlTgzHtytGtF1L7n6diC+JCXR7SpTbm3TsZVFVIwgN77jujhedQpm3S1BCGnk/
WMfcRM4H1lBE7h9uzcd6zGOhZp86T35rQb0KotGT9A/A4kVfpUb31bvN1reHxODKITckNQAHbj2G
d9ks+9XRktoBroBPekb9ZH1XQf92v4o/jqXDoJ7NctyITdOyb/Ax73ql5noYl8Lh5sCpxCq2LO7k
EJnuADas/lbMf22KU3FuX++hjS4LqUuf3HWbWT1NntIcDppn7Ld4J2FQkhmzYN+uZSmgFQkhuYFd
NGh1JgO8cJvYQEtkdq3rYMeCitZtYsHj6ta9ziQODyansvc+wJ42xpSLYFUeaDAhRjrRBAV6vI/a
1cZhEJ5ZWPYVYFmeX0hKHcxe3+TIHq/Q/5V4mItGaxG+cUsvlLDwFGE/wHiCQ+CXBz8SHzEa2+nj
eAEQBPgGL8GrN/YZgTDNXY//1DhUFW+Iievbn0shxSvCHjlgLnyK4/cXAKjp1xwoSZmsZ/j4IaQq
03eIG6DqkUEV7uawzniISBkeoP9WV+7Cu6ZrkQOjgDbcvor3Ib46fxtdb/zaPt/gmUk7VvW6ayH2
CNoL7VJOCyELbHKPQTSF944aMJg4MD4DSKafiAhCulznPhdjTAb52/lj1VLcw6yTCS9jP7Igzefn
Adi0LCZJoun1tRNek0xDhNRhVYIA8V0ucTMDXne4LI1oVsqax0rx0Z1m/obT+wvyqceAbbIuvHRI
AiH+bBEqOTTIBIS24HrbkEGXSunjUyWFOQNqk9USZxfEeiKXi8pDIq4t5mXTQzdjHXY6W6klfKcm
ULUsA+IWDbzHhOxf16R2mIPdJlvySnefuD+nuq6PMvohip6xG28KLTYSCTmwBGNiq3g7rfoYSYBF
RDrbUk6zSifekBVJgqY8yjGKvXcpeBnZLvOyn85YuZO++ryur/Oa/vQlSEZq1+bat+Ez/vDW6xuZ
Y6Mlh3B+5jC74QINJeAmxi56bvvQ2y5il8stOUqoMlYkH5j02Xkdxidb39b9UTpBCaXOEBwiEvPR
nlIXn4IFHiEw6krkRmadzW5cdnbxpT1nAdRzBm0HDS4BjdSZfrvRWvYHTrcwoBi6WJk2UEymrQdn
pFeBWRMfosswe9F7T/HKbN34qtS5UeRd6kJZvEf44Lj/5VRd7Xko8SnIO7VtzCVnrLQD5kpYiat8
5y0ju3/DDnsEWd5yhcLD0uFjnpOqxuPEIhkpDY3LL30oM6efvtrIjpJzX4qODcleXwiZLNrM7iuI
6tM6i/nWpHcxqxhybDgDn5e7GGHZFLjTJWXgu4HD2cistv+GSFg5BEDGGsqUV7Qaf0CCCIO0RMxh
YIo7mjMIxlFS62Xxr7+zz6oixcqkJPng7QWyPQ6ndjJr/OS8RbcjB0kMBPsyhgl/uItrMaga6esP
kWnYjLG6nCMDSLnIffnDAhqjj1BYjXKrVCNMfvVnQ0DAFec5L604Cg40cxNKImeJsgpMXKR2M3Ty
0Kt4F4R+IJL6WRmcG7J8tNm+h515kh7XXm8GbRjc9k5/eykb9M5YwGpGWzMswPnvTnVCo44v+Mf1
de5vEwKlHGtatLzEdrSWtT67shtWiO7NOqUQWcRxmphNVfmiB1qgzxR21QIdxpPQ4MX591uqtGLw
7Wp6QlUIydA2HzTTdo1JuTy6ycp3cVnZLh36vSYLy4Fip47JdRRlGCJIt2KeyZyAYE+9Zh7x/v3x
2DCZs+HWTbEXGDmysnEpr4OZ8V5RVKl/u+JjA6T0yZIVNhisvnqNJtLj87OAhmJeRXMK6jlbRB+g
r0f50vAdarYD2WdlGIiTttH+x25Nuld9Wc4vkZYzflmWrSPPgPAp5tvZb/4s+qPIy88BMjAyDNmu
OoZt3fayhrlGrJsj3i9Oads9XQj+9cOJZZorOiKa8z+p0OdljEue86UUDLUD5zJZATxweAFoch2r
IuhQQqrU/oUk1FgEWvbWLmXrlYe5qX/OnLxwMOlc+0w5EiCGOSvlqsdvDQSltoJLk7jD83LzXW8+
lHPuoEa3nKMJCZSLPoThqIN36qV5Q1M1rgGokozGyBwP8Z7v+Kr7Sibifxqe/WIqZ7Kz2un2TIAN
+spPtyYQt99BYDInWZtDuzbJg/AedYSPL4uhHIdmMLdrXGuW3GaHCD3+JBZaE1FlI/s40VbL4oBg
mfT2NPzYc+cBCJb1tK2ksea2qGcegBlW71WfsiKnAIBFuACUn4HTsx4gvRIcGLZBkDzaKQX9DXAR
OI+DUiwxcaSmteokaaOaFbEwrKwBg9xAZjJ/Lb8y17+75BNKwid6UJCqCbHtqIdbMAbkkEC8nPoH
jF3YOPWVhWiZ+cMi7vdDQh6yh6OfEeOyKwXw00reH1mrGDv6Df4PjS5yXlsTsT6dWH64Wp3HmOPH
PwgKvPdBeIJq/CD/vIJtVSjur1mUlutfU1+DyIJncWMg+5B/LeeRL3lvjISwt+pLFP4vqBUS8HYQ
KfNMYU6ZrmdWoLVs9Nn4lpUKaCf/hwofgthXfW49bFt/WMepa+r+Rf8RcJ6KnTDlS+8HXepMlOWm
Wxqc2i9V9HycJ8kQvvUlDxqbdAxUS3cCxwX8knyjdftMSxM8AHusxfjAB0R2HEgPoK0CNDAvVh94
gEn2zT+3DaNByWvDdN2HiEwbFW2ETwGGt5ObSiwj1GOB1+KJoQCLBGhkrnNNCxoEJy2Q/QV1Rdlh
y7RlJvE24eqkJRA91A0EJ85QiIuf5l9tnpBqplVaETK5oFWlDHUMq4zpwiCUlJuoaZmzahGkyWIN
3NQ74l2omaih5n45hqwjGJxqJs1VhIaH6mkrrBq7U77XPp+2laotl/aaGYlu1dPlAI3wvGBr2B4d
1jdxJ6N2cqfzE+8JYpBM+JARPrxmpm2DRl/5IJ5hxEpvfdOSdOYDgMUBr94yM79VQD0QKYfRyu7F
uZoKvA0WItzNN6fmiwvpN4Tpgw3VIaX2h7issfd3uBHt10Qjvpp9ua5/s5I8gmk3pHeDo4JPhfLv
CCoI34680XYjNtLClzwkpFvKf9GNITazl7eUEFBdx+BXoReAxF+rnqy44ARI1FN2s9Sa2Fp/GZZO
gSOhzz2+diRfkJxDx4tZaFgXz+gs4zLchEMJrrXbSxF7FrHZD0BRNVy9AmZOgJWzUHo9E7hoZD7I
MbQ3UcdKu+nx6TvI476t8TDgK0WoUVKGhMFdX27Pwor1r/ErgpdDi01/v0p30ylui2hTgJkdx7x+
pE/3yZlHlqVY4UhHiyg7yHaAtAH0kt3IbYgcBJuIqjxmr6hHYaSCGVFYICQmHvyB9fwjwMBuz6YG
DYBwzbys4IwqtND+0Q5W1umTEvuuzAn7WJAsnAXF8vTuKZu1H8RnoGUmBFE4jFgSrXUzSHgR+TQ9
lsrPrVvBaVsfQ6CfSa+ww2vXTjWa7Z5mIW3uCzY02UZSGba6h0kbnpALrkbR3/Z6+OpDdnYqOTI7
lueuReuXBTy6gLJ9u5BJlgZJC206MXZLDB+TcFqYNdlFbvKCVdkC7VRUVFjur8QbpBCFBHog4Iww
BmIrFnyyP/quJoQGjGjbdheKvzHMR7zCzXrlJLAkf2xm37PDgt53jbrBNKUo6yQ28CbQz3WV4tWU
pQBWcvqjKml10rYhXkJzm+lxcTq+Cjp3zXq8HP8kY1I3CE04sfpF4D7Oenv88EIhtR50byHNToap
aUEW4WFp0IX2TEhfZIjncwaPHgh2uQXDt8YeoRK/KPn86DDnbpEfxdHID6M1VEmVUkFRfXLwLWUu
Lse1pzWrlrWP7hVmtVcQl28glu2tqwq755e6FqqWd3z4dvfnQP8p+rbcnpBvUmrUffgTx86ivOjo
Z3Mi7wKIt2bFjC5P+O+veKupP8aiZlUyMdYeOgMh/x8uB5UgEF2oOHhtadsy4a/e+5U5mBUHe8Gv
UtoBeSkUKgOH6AVXT15trUibGFY1k0PS6unpA7V1KhzMlApmonnBSFXWqQIxaYAP4KW/c9CTmHWm
k/sXFvRs4XWmZNCoAhxcAEcxPzutNIiH+BrLYp185URD9uH/vHN3vyVA6c6v6e1dwddO2sWl9Ese
ZLdHuOtZAJrhbJy3eUjulyzjMuPigjt27W70WNH2gMNzSWx+icNYO5Odqj6Fxw0/uG6oN+EsGMqC
uU4FC9VfaiQ5iaewJNwz6AX/m24DjSDV5pCf7QbUssmdIph0p9EQUMjZBXFrPLE2Ow4blHj/fisu
ccljU56dkfARbDWuR/kjCW9Pkha7SESjz3rotF9+5Ksqrw1itO4vqqa36aAH++NbQJNoXKAO92Pi
U1+4Z6SaTArNrK3Xw4cb4LjlCHodm9RtwCb7tmejS47KBr2qAajWjGgn9RM7Ug79Ml7ehPCPanz0
jb8ptCIZNgxibV01LuRO9jujwAZvb/lrScBg0iBrdKfzHeytp9elRFsTrDyiapFqt/5mBA7RwNbm
AwXUzIBe0DUvNLStQL1IIVQkZ621EpUxh6bcxtsqjiPO68sCQPllbQphqtctFskLonRpeCMKv8Zi
2Q0Sk6tin06x3WCpoczA0pu89kcNFayGZB+rVZ3S2r5/Xy2NouEcrTkZ5FyKEQYK+17YfbSzLzzH
qmviAqCzPs9vmMtAp4tlyUQlZlmq6zF9r3C4oFWk7tjoa4JJP8mL+/7Tcgfc0dys4vYj6kl/mof2
yoLGavtm6O6PYJW4qciv3Q9jh3Ic/OEp1JyWOITRXhdX4wT0zwe17ztrrk4O5WRZwCHxZmDc8jrO
OG187QntolrVdUiQ4T+tlU4nMgdBNooEYaIIu0wonf2NbEdxo+urUsBxHcgKzwkSWWlyAs0yHM1j
YBdmcGD+cnh1NPtpUQd5D+6jdfn7R7gG8nec0+MqDTFbqNzfm7p9mA3v6lMcHfKa9/BrYO0CwYeh
y2jidnlH3bR/PlUO8nuKGu0vFdduw8h5zEtYe81I/axssv2LeTz2Nj/8FqdwyJIpYq5OELGNZieG
1Iekb4mupK5v31x6cwxtLd4i0kmTtDCsjFH3eyvlNOdESvK1mKHv0BjpQLwEtFCBH+cv9Cr6HlDa
FMKoye5QUAC168arF22sz7oUeC/arnv1ft23LPtSmHOM9ERiOEVkbxilX5lS+pWqOOO4UVgmoVS2
r15XQX4OFwo9SuJKZdj7G7Qqg0IRAaODhfRUqcLFPP/gcodP3uZ2IF62AHCsSMgJUYx09kwSv68j
YP4Vbb2yiUAz7OdlBCeGLCYZDIH4eSKEGwD9DglktEB++D4JvHFCq5p7XvQfbrxIiv+qJvKHPib5
RIoU3tDU8M6OnxGydaVi4nEcRdcVfhgsz+yyqdri2lRscxvsHt+x8nFGokBJKEselh66kSQBwoF6
9fsyrSLOZnX7es9orWbvd6LqiUkEzxwi2VzZXj1It89EWjoRArWwxVLdCdHsz2q53DDs2mqHPLzK
pieen89LTLo0R0JGC+EXx8UKfYx/YWi+9aaaeFE3UdK3RtusuohqYwMVpZHdiGK0jKR372W/TPJv
aG6b5SgUp1hZZu0muH4IcoEToAN/4w1bz44waQFSKHBAYHiKXhKAeRttdVeVgHcxBqm7WcI3LmU2
+A48S3N/rKmLjcdcA1TVfQBsMCIPMEWovL5zzEkKqczG8MK0rzqKsBUONCjOzIslVQlJKMzd40+A
dQekeBhkmgN3wzidOVrKOALxt7M8mvndTc79rXqMsLqlfvh0yJC+mPRUN/0l6iF6K8vT9GjcXWD2
vHsLehHw+fV1J22/IbVxmpBS5dX6vRnmgdR70f+hxveoOLOEqllCtaKNbWVc/a+lPrO6IkJbm054
uCir58qDHAJ2OyRRoLirMF3F615AFVDU4P7MXwZLk/o+fTEWclfYnDXuW5fqvGHEA8Ms4NB25MAa
VsNm5yJzk0ib7gl1/Js22JKOZOC6HsrDPB4eWs72/rmK0d5IXD6OPbDH/HuIn0K94QCa8HplEUcb
7tRrsoxJGVaNrrZpcRaiIN3JOyQoLr0aTFIOVWLW+6BUQTBy7xhtEaJBlLqfd0d818rnYo2s+oVc
8QgeqjIQLqxjHSFyUMkimig8cZROo72lqd6dIFpeH8zrvzRm6QkAHE9dwaGRJr0hYEam7M/JaieN
XtNWmWYv/f7Oc5T6R8XXSs14PMTTOMMwUwXqROWUCZYazdUqMNUuw/i1uFQ9uJ0dnm+QgKSQwBbV
FHFQ79gSfbG8p1q9M3/Qq3+s1o10xcLz2movAwQxrkWBoLGg6Z1ywG4gcuUIFULTUhpBF2u2WGP4
238Hz+4pLPBvMa+E7qj/TzojNkG9BBCN/Epq/QfZ5M7YtKiYk2OAZgwkNo5OVfcpOhWgUNuul+37
8iz9Uy+HJB0Q2hEBZHaU9xx5aVmTxI64Oz/3Ja9O/8yxFDkhyMxDCTNVUKRbgnJb+MdXmUQXC0v1
JkK59pL3zb9KdXMBomjHR9ft2bEsbJVtCzuMoI5Qgqe5d08Fg7jPeb59QPOsE56aIujVID2XbJv2
EmK3aBPFwrUNu2/k3j5cUKqluApXdNRJt7Vj/n1fBHhbNvKsI7hls5XtiHLWZZNB9GSqRvyBSfNx
Aie9fr1Dyl7f3QefAbPJ/m2lOs/0b+GxclLKrKiJhnKR2slZqRkWavLSS87gRaCWAi6Ydorlnazn
kW7SEXg590duuT/eoqQ90a2eRrbmcokcgeHeLhhrKcXSS8+3hsHYctOwifsBq6AKrmkixyti0WkX
jkvIXFrGueE/1N0iUA9340juiiOgao4vUdAP0X1QX+bGecKdgFbb8wPl8uzdvaKjff1rwLJpGROl
nOHxeGd24nAsRa2BBAXfpPAFxOzjniXPmrX8IS8BU0GEuct2mPVjmW0A/YVlC6cR+DuOjVsoN58J
oXuXZ1Q+n4s9ATNod7DXNtkvAhvfuoj+1m0y30un7a50HfFGw/p+GH4W5st4T+5ciNhPqggcmYJL
xPyO/Lrt5AgaAsxAn1zzQOI+CJ0D8bWFSwnaDZuMecdHJntxW2tHdhT6ldfGMMEejNcZHxH9aftk
kWRVvsBgG3MWRAX34iVdXO7wIq58fSJA+83cH8D6YIgpNMtid/nGE1jkcaVcB0s8YktF1EOZ8gsO
j01xZtMGokxJjJgauA30zBz7YKD8J8GW53vxQJ1lS8AycHqShbVb0cjFHrBd2BoGw030E3zF33Ui
llWHl0CpSkpXRR7498qkBBMHJHEMTzA0VDFKJjq0CbnbKbKKb4EGYvb7i+y9S28rbvtRTXKtvEw1
PsGnxtuzgzF432ueo8iOqm+5da0gUFcTOmWCrxrsyXQh3j6U9wWLTvDF8Hc+pFIrNEnn0hL575mk
YcAiglSIcs3Ep6Mxj7eFCo7t7Qfaje0eMqY36bWi84p3skC4WoTYn6Wiit94MUuRFKntqkP5fLje
E4DnRgUONdUYfH6ac/wmj+SFSfKNsybx7kF7WS/EyhlN6jvq/aqqTjDgVN0pBUrDsncT86/L/Oz4
ncn6PHV2/lYkWroWhWMXinFOoBZvR7melvRWFWIuUFCujuc3g7lCSWnpvP2g2vDmYfGLW8jPjzPT
cUgAb++Cvm66HJ0mReSUuSlr7gH+0Wz8BXRmnPSm5cHDlxr1RVPu5lAqP7l/jM5+mSf/sp81vhus
B4g2zJ6WoVRax+CljJTlD/JBRJh5g5n/pYtCWVX3kV/HDevr/5FXxRHQSGVMm/sdLbHy/Y8DhKrR
rHvBm64wtvp3P/048ednZpPVqWsMk5on1/LePE61n3EJK86XnRCIvLL+AOP5byA5P+RROdDDv14T
oCGs++YYWE/rwqecqwZChwgkjqJzrnVpp6dNd8Kkas+h1k+wLxfWnm7SUP33k4ta95mFN4ybFOMB
Bjj5Veh2tnfQt5N5RX9ybKAqqpDnn6xh1oVubp3wFfOjB1E6naZRViYRuxpaYKS8rTfEWHELhF1m
EbeBOqWMk9CPGhai6aVGP+VVk6PBXN2hGB484U7koYqJA+uSAu3f+Zat1kpE5LwnDMrK+eRXguLJ
2zvYVtqM6siGreBzNJzg0hkOhXueF20gNRRx8bs4eyGu9gqPvSjfwsjJ0M57Sc+L86Ily2H97INi
k9UR8Qysmv3wQcP0w6xpAko71w6tIhG9sSXg8zGIV3gY6eTgHWG5G1BQLAcrDU9CqUCz9/nD1P5/
FtQTZX2PdqUgILFKCirdYcXw3kqtakH0L5QCOENsLYoyYDtLFwXmpq4h/fxv854vbdare4DZ8WSM
UkVmel1rBBWNSnXpywBGSXIOGqYBMU0YAogche8Lai2b92FeAZ3/J9YFdO4FuP8McmN3iN1wtLeF
hM0OZe7VQSaM4MW7mDBooVFzK87kSfpV0zHLSkPrHAYPJzqXC6U+WhkoHEcrBDFdghojYdXOre/Z
BRIcinjMGBtWBhFNLBBBaOrbOHMb196TLt9JCzNvqgw5xWVwTJ2Ay9d6OS2KAZ+82U99/XfoD158
AxyvSaDho5GjtDNf+oFxkGolaGEfZQA4N4cWbHvvNLQCdZ63FrPnyIhvaH70WAwr1dZ3ZAGpnE3D
Ed9H0FQa8PN7Y2R4dlvTm36Xk1qi5+xOk4aXcz1nJ0hOveCx224Efa519fuRJA9l63JRgpMPtFaY
mXgFsPqHlRRh9uG2MuqJtCwcIC1v2Ol5JP1SnwknlXU3J9/0a4cdUqJmlPSKM8jBYADd3R5smpe5
WrQKOP7eStoPqXQLDWV8XrW+3yMGqrWbQpkOWa4TFV9zK7YvDR6mZMY7wfwxctYmwiSqzcmKvmZP
J0PkXLSw51bwzGsY8XGU193R7vGzD+4QI5USMv6n4O6gF4V4exOztZD6ZkanLDEOzynzLzRyNvji
oCoVIGj730j1vkwz+Rlg6G4ts5GSDUd1maYcaQ7qdSH7hGKtD3CDitIlAL66sEew3Qsl5puBF0GX
ZLz4RWmU5ODl/8mVxPjKhbPTOT57ogmI/u63uiR6BLbd9HrAwuBmdFr/q42aBRDu2BNcMMXO8iOK
JTNnPrKxbrJPPBAkNXqL+PY3hhKhkyqEoBc24doWp5+loExEHD+hE6+gtiQtUaC6bNIjNRshJXgd
xjnqKejBLAMAHS6B+EHDgD/mVGnPpu9QFRgQqouXGW8EUY6nN3i0ifMmnY/4tzGwXcfDXBEuqoYa
2YAezS02EqNabnCcmzFg1SCTvWcB48nR5Ts89vfa02prPOJd8nJXh+2Kyod+SASFhSgdBLJGkocu
K19eyGuLxSXxwq5u7ewH5Ib3PqVMyQFL6gup+zUSZUdeUmI0UlTO3csQ01dYMuIBcy6QiEINX9x4
WM3lq4wPtFsSbsnBcpZombb1X0ZJls84DEdhblWZglnKd4EWFogRhvPwu7yGBrqzCokkAxM/Ez5d
P0UOKDNIiXLsKQ/O8gsrwcE6Uvfv1OECIifHZ5OTJiyaXI7B0vuVCBflc8pK5kgqqZCK8lT3MKju
/lB09lRJgCY54inwiZ4q/8oKZDbWgZxMXzwFNZ/Y7YBsuWnVW1+1y91DQLCSs28LLZ2JTERSlESQ
FBcVv0hhTBGVrVU+7yqxxqO7M7W1WxFBk1ZTqxIipry/fnp95PakxOP/KkIeJvVEAkJxvrY7hLUB
P6XjC2pP1KdxsGKBPBIVCzI5R+gMNXrMw9JM2WNzRglNjBucr35FvQzdiqamEpa6xlnXc4xjL5MW
VsiuY1H4Kd6XIuMsuEPM1KhQHmhZGKnDXf9DG0uyw53ieZi7JkJZr5IzrJA9EZGJDy53ip7wvDeA
sDxzqs8AkIABO3TIleJ2vxf8m2Lc9ZI7v1ebBpEPz686dUT2WhuPdXos/bHkzsYoJWsKOxqRClsP
QsUJUzb9i3OCLq6zAWHk1HxtSiZSRgZCKEm6DKXuXojI1b5YE0kcjAmd9btRzvraYQ0CF4xYjz/B
izTQZ7AdsEQjFbBwRtVCqL4JfZe8sXq2s6Tf2JgP/YL05x+iGp/23BSkB1nY7WPYRZ/4TqBNIAnG
DDlr48dPI/BTH324l6nVGx+eDuWYU6lAKuDwA0ycMLy3NwpkozJ+HsqBDfVQMTErwzHbXK4hj/Cz
+ywox6/79Jp/FgNDqSKORjnuzRqQhiYtQoEryHrzKHzYK2c4dx2oe2IZZ6z8FPZ21tLbJ9GX8Ze0
O3a24o+ngf4XtHdElVXXVsFPoeK0oCaUCK3ScnX8DLJrm4lPb3Hv2kLj9JvPSzMsLc5Vy1gZq9WY
ewYcj+Wj8XFUECw6SvSkFtFRqEwVsenkMRilo5VFVFgfVLvWH41FuMWY1BZDmYUN+iqwCy2x5vx3
70DimNDxAABvK59+svEz7Br4/8+QqQLJc6+/nKHBgNxa3mjGcBGBpyl0oRGJQWlQhliIaZRqv3eC
m7EZNM9TXPWaC/CB0//a0DNa/tPes7Lgel/eKTV/Sj1BZR00B4ZtBA1S+BVOsjCctCwCFPeFfr8G
mZj+PkTa3nLrwBbaHkcJcSidCNUS0o6Hh3wHJs0zqaNBUdnMuAosRxfEHHW9F0J8mDRq+FC/izGh
gkkfcDkPQNl+1OHIpp/vAX9NPWSE5N6T+OlJGSI6l9BpYBmhXzcAc3uXoAXtOLa2v+yfhC8kBw8w
012AG/npkfWXvdkMWRwkvV+cnFaVPMN6ZZbuKJC6HRfsL73CBGnRgBk9lVAaRahkXrTJGt1IyY3s
rwa6cqRs6gq04NUyK+VcK1cqQGBQF/HefxqFff8Gt8n/scXjCzFp+gYfyYDj/DHHkOuRXMW32tgG
dgp/PGy9zNwF5kTcR95BGYs4QnV8ZXvH7ZIzGdd5rIMpoifjsNFxUkEcdvtxW6iFDmTEGr/UKFrD
9Qhif2wA+CkB4paFCQsexOGshsSL7R+Sale/40r0F1/CCnf/S+VJWxlOaAW3QurYzrY3oFBu/nVs
fmXpehy19ufCDZ1ZUPODDb8ecMak5tSjN87oTyhYM5lpbGMyWiL3FpOVcsV+Cw0jrD+PS1S9ZVE2
z4sol/wNxmIYNTyCiumahGB+6P4eEjQSDJUYWuVqCjBJvzCyfsk5TWsKiY3o+cPhIgyzpGFrjmOC
cxHzShRpGg74m9ZQ7TKme8rQfxpIXBWPJJka3T5BqYdHH7fqMGgtlTbhTIz9XZxlF1kxmwdWZvJ+
JsroBq7idthix5EVpN6zyymRKLRsVwh2MQBXd0N+bcOPgViU2yKyabIwvFVC8aWOAJR6V4msY/TN
IohhpER2XWewiI7bFc1dcrgdLcjinFpVWoZQSZEkp5w4PLvTYERMlXp+4ETL+4bQDie3BBCi9s35
DGJsCQ7e5TY1R/bxSUdxBE2Qmp9mQCJnSfbE6eBMmVyfV5uFAtrUJhnYWQkuTGz0lZfbcDcZS/uE
xHT/lJECHzlpYlY7f5xu8apbBuX/tHs6oNAKJU1C+ssecvEF5Yufm40LFhYHi0YIG/JRb468Um5k
I7Tv1W85HhYwg+EXyxtdfqs5sB3comb4zRaTOmjq0bw9XirmgJxSA+hYqI4b2ygHLgv8LYiQj5OY
F3YkOj4IDUErZrFKyx5PdA9LgGcWhXU+vR2TqW7LzxGiL22mH+Wta82Z1/TiCNQK+vI+p+ZA+L+y
bB7TskKvfr6wEhw1Rb+eijB6oNhtScUfnUnOY3zFqyoWbXQp0/Y/yD9Ozq1FiqtrAh44ihGDckhy
TWNSLFUuPORusOWuEfWBtKDvJ3DQElVUmYPXiGSCK25+OgrnCCwPHOsIFp2hSmMpO5LUKYCUDWnM
gzihoqdMUQlHJcKhXDf3VeiGlAOXh1gynWCclJ/7hSina1ztQkfwSIzNanJL2r6NFOx9hGolZQXt
ZpICHnYYHnlTlOS031uPtz4Dt8+c9cVl1+WdvN32lteFle6JMHB7UcbAWLmt2x6pXlV9bl359iFd
1AtXCg4y4dYBoceS17L5HZtPZddC7T4xMofggyQ/CEAe9t2auh1qSCWEZCREAEKA+8yK0XXaCGbx
89iGUBu+qhESvtzdQxuyAtHKl9qwiqaSxy8WSAo6m9RHdSS99Rx/cCVNFn+TODf0VDEelYp1tOWO
BjQI4UUCf/5fyjNScB+bVVKRE31bo6zCzJKLq69gjxcWtNN00jUtP2mYWmaf2CmBKK6qwexBlqsp
GHwy3vx2DlGKlR9rJttwgaaeW0MlbvHDUjbtQmLnEMdUDaxlLKCU+W9bC4aix8XGMUA8rsIZ4Q2O
B1XbHfr5SBviA8ARiPMVUWlz0B2S4m7ycQGFQUaXKWj5ra9p/TAq1yFHwYA+wvuqH+UPMLMRJHrI
PFo/I2O4MYoNW0tl60F3CljfOG6AJ5KX8CfkvyjjrIxJK/KWOBIiyGNpSh/Kg12lLrsp/unT/FKY
o/1h8YQ8YGoPPwrYBrFjSbzXJo/B5Gzt59VxQ6QfWxi0DIDn+zMHy0G3Y0TGi3BuVjp9KDcpgktd
lsEAXRpPBcrZVRISuuaMgtQV6ZgcwFydkqeFm2u2RJlHo9nA7TYNfByh0zxReHWPmYP/IInJJzw5
T5ZSsouX+EJa/+O4vor9jv1ZW796n1zEDRLdVvIs30R99VhIUo1PsNUFTIKn0L2Dk+rf2gCf0Pal
ELIb5D1DumW8hgsBUsojvyfd/RLjPS1GtIuLjMeMAURl2IcR9FxgFZNW6FpX1zZbsRar/WNKxpNH
bq1Hlxnnbg5yELpp5uvZANADznhuDwGrDNQn/BcdmL2havEA0UNLX1E1wwaf2lQWzRuzDw4+Ixai
AF3pMZI+qKLSBrXoBRhl0p68xhXZs9gsYChynu6/VmL458sR2Bzq68Wv7+ln6pcMHuaoSlMDtbQi
OgYPqN3bCiOVtjCQF8F3v1hbve6XHI78jlB9lhfIs/MOhZUq4EAI+/ktQr1ItmWyLyVv9KqCLIAK
/7s2TSV0iK/j2r8/thIms09jZMaTkqhU+PbwHIx2SLalnODR2s88NzfwEOJLtoZLXUHXvc41d/Kr
ixYZxf+gVDULrM0FPJnyTFcpPRBeHYrVwVWrXb7fIlq04R408ZlQCsWPWLHJZXQq5hMd1WwvyDAW
p+dHHr+/thoKL03qipiBQ4Q+LZ1R5WBYCu3WC+Hay2hkV8cacMrNSnEARW8rj4SBODpTxbxkJnDU
us2SlDK1WMJ2CvNpp5daaMv7p7mziAcKgtSTOl894ek9ACJIK3fOzPTZL27gtPpJ09lPx1m1jeQL
GA+8Ugz7mqGwwsl28xIimwzQ2xu8j2lP1ElVdqWw5xZ73b2zjFrmGeRHDOsytwbCb+otjtXzK34Y
RReW39ECDLaY1QuPSNQA5Pgfw/ylZzGEhjtb4Xsn3hqorKEwDSQk8xw1XVk/fmfipw9sl+vxPHde
CBywHykboxuq1TfmDqb5VQN4S/eKhfLo/UAm4xlY2N4+RKIRnYPGtVujsYRxpRQhD2lGnfstxMR0
4qqB92w4smZAY9094SpKAyUipse23WrTtqWAHeUHiKrqY82NaOchgmuq9Ii1nCALjFhLnP4Qb6Pe
RuB38Z/0y6AZryyfbVB7PP0yC406tTl/XuIwU5aRNopXcpo6VjwvNNZLQwY6K6Q0JFzxafYq9vOS
6NuuaSqnjB87q0G24tYruxRDOhT8dcHeAozRLGsoQUocneyIYh0lqGQxkuVbNkD7IbW/zx/ofeWh
oritW1cb0v9t52DkccqFnrA7pMX+5AB19G4Kb8x3bsJ0LU0k9oNr+ZYlKjkjXmDBxFYQ8UPTDekN
zIlvHUJ1zlWLqNxqXvxl0xJ++6uhL4+PcVW66h6G7xCLds81QmsDD443hjLAe4SceBH93DA9UbfF
2xWJlPm8JXfC5fNYAtoP37PQge2VTjo6nkjYtHOm9imb+fPWWAeKTjcQdlna+poYGtV4Di4sicge
QZ9Dq3Om3YAr+Ui4JrsAMAKjHlTTPdF4nSYCLHXi7GuKCJsQ0D3eXzByhJlhV9NJpp6mw9+hmn8C
GQlmkHj2GBEIaCM/EiNSXOky38RCN5XYjtJIHeGMFXdCtun4URrVt4993oANM1K+8n2U+kuhAGJb
cSA/2HLz5/duDqBOR5OTMJsD4kiQcFfqqX3nA/J9NqifiwUP2IQ82tR75wMkRpunsafsm3xbgPgo
fyaxDGG6YSaxrWfvM+wXPs2yzwJmOTjvBXhXZiSLbM0IS2BFy16tGD7/KeouiLUZ3iWMEOk3tfW6
s90TiZ9GOkA7XriAU40wb3GLgomSXpJyA7fHovHgXjQ4ZdmQcI+zZ2ehEW3ZJDTVgmu85UiF+PcX
cUkBtisEsVG84pXBH0hmYM4zRgok7jABUWuQLoZ7gdPuyWP28AZMtm2fsjkx+G/HM9ksBJVv4vhG
d1gLiKbwrrzw93n4son1p66R5pa6P2PMxPCNZew4SXPLowvD+NMswa8q258eJxiRLhDrWkL6iaFe
/DLgQ3VEC2PAfZN39KOhb4hs5hDg3rOfm2PCFhki+GzSZlIUcSNVKmbYkybWdEV1RkYEF6smmHA7
IN4pecJuu86v//ox/QgibwQnTrbkzHpJzlV8e6lpAu5a7At0TA1RvngpTWRgdb7R5/GlYkfExUCY
eEyf9qfEKuFX2WbztSPm3RTDxUiLiFbLSIlyXAO0bgKBgLHy0qh4YK0DSm4AsRogXnkdidKCCjZZ
HlkYdiyOgbsfQny0ylqPMTkgCMouZusyja++SdAMBh9oqWvyK0J3FDQ3JdJdpOw7qkuqwVX2ziBl
oVMG9Pk7PgqAOZQbDBV9YKNkrOqX9VYN2gkQFfW/xt9qxnzaRD2kL1Us8qtrgaLMJOYrnBm/NUqI
Fm0z2SmpQ1/CntOR8kFghJhbCtT6vozlEe6w+RPoRxJeTcF8xOFUxiEIWqLWHb2FFZ6b0l5Ajnxq
+SlBY/2fw4qpHbhw9ePOHxcgnagTBFIcklPRzXTUBlUhX2ewLxk+GM9ajQARJv3Bgk+7bAG+xEZ4
11iMSjd+LusmBgiKXDlbG6hYEnh7/bMCgXGQFw9ygvT7nqoyZro3fxHJ8IthKzy0WZy3XOdxHy4W
cj/IvM+tHatBqWAywFpFLNdA+WK6UTh7lo9aQ/BaYw5WZM0tskNFAeyAVUdgsX2bAENKivvDpT6r
4As8QF2I+SHCJdBNV2iVK008XIzf9WyOcJjQZT3uy0gSAQy12crCa33ROWvGKzxhF7DmWvGgM/1Y
pyI2hku4m4Z27e8XL1axJs7EV9+2C53CHfs/yHD+Rx1S/vCp5ZUlE/U2DoD2mz1FeEtO1AHmjw87
rv+Raii7FIu7M3WrMhkU2OAy8RugkMObpCUZSrqc9xx7RPYUhj+aH5WwUg+wTKLAt6cvMpMNA9mz
9l3SwmYPyyjkmbZ8JEXfBjWa6qnPB/eXEvYaBHQsDp+WXz13Peu9kp20v4kZMUHNdGddraytT1WR
wSqoxcE1znpZo7TitOdP+srPAw751nAGxKf/C29rRAuJHWRLtAGF8Gv9ZQZB8HTsoktIfI5Yw1zn
f1x3DTnmMDyed+R6UD3fvCzXe30m4K1dJqtuBaMwGPHwt3wG2RHel8EhjffyhsBFozRqh7QdfR+a
EVnRQ/7Ztq+UCOBP7mRxu0LQX392uARRNC0aI1D+rvOQCmm8znpLUeWlLknc/r6TaJCRGBvUZjAB
iZxqyi+rfaFXBscVENJT+EIbXXGCgpwJ+XxqIxNEwSyKF+LbV22bWHUfWEBDyJPFZfu5CDHR/qMw
cOy27S8nTFzqlIgvL/dC3T0pK/CA60n0r5EXz9MnQk83zudALyPivAkySe3E3WnXZbzg+kqg5/o5
sGe82H/hULwJtcvHJjefGUQwUSSIWq30zD+8bY/aBp1wRuhnA+p4lEEQiLqAaEzG7rN/gYcaVNDn
BesP2iYmXzOY+zQbCfHL/tPHQgjGbGsHsN30p3IFq6DQT63SIKFaVd6I/tfGKIQEyOKRg7UaZkv2
7rgx0eBZ5QLwIwzDdVqZcBzn+AZLLXYPGt6FfpjBIYs+1Hpsvg3GZEesyGkjoPaEAB4se2yylGwD
ptmh4aLYkalzYXoQxg6kSwNcgYWwvwdf3k5OMvpI5edEuUuBg1dZaW0IUF5ILZ0jYIBmBi7zAyNr
B73CWizksMz2XQF+69fxK58KlA6PRJBi7BzrBSO1dk6gTIj/gFrA9/5sHnhOuniqULckEq/dhK2u
qq8/vW+zBTz8x+MNVBDmYlXW107TSgdAnzBu7GQ/Y/drQaUU2QIzdKEECAdU+zi3ycgiIiolBzSb
Ud9QS30RIr8o5N2p41SG9oB0odL/E3XOdBjDiMGw/NQOd9joCSfTGl5ym2mQBIvVIkBVkKL4fCmX
gcpzIzTcl7uoFTwYctDloL45wy/YAfNud4BjLnoxMtSTgXuP6nTz8YDFlollwFHl/5NETyiIX1Zf
d9da8Bj+JUETclz9WmmK8Cg81Dv9ehOEMiuWz2+Org6oukb6zZN8ESOhDuT00I0e4tGOJ3L9CxGa
78wT2kY8yzCvjmDubxwSd1n3AET43T92QkxK7WV3xrVELhSS0CBGNtugK3P9VcdHBBJJS69JG5kp
OKJMo0rwZHAMN7tN9sRjAqfB0QdXF1b3P75yC60svyedAgfdVXdzAKyjo3TnT6ZnCcjDmHcBrnGB
QeezS+/g0sUC9n+ImB2aZLHslZtLlgz9wmFDa6nMl5R/dy+suflPcQCvdTyzLBAKntZ+xsqzJrmP
hiXYIPqM/QRMD2t62EzapGCz0cbJIQsgeiq+MA0ZQk0qOGOg5e4ku3q6/m9GI3dDnbm60rlAi7oW
fgJHqgeGBw/I6S5iKndKzSlbsBDiYIZSyzTxK24JzrDBPzrQUutMmo/vNGYjuBDXR1VCqOXU+VnW
zar3loAEtHmrIeVIOdQfO3yM+YvMwIAqrLeqQMztA//aRzHpoTAVNOgWwTUH653Dvwa5nEs+T9za
ka10GZoz8b2/fXVzWcDUwTMKr9D1YdHkIZ3P3fowdugXmWOYApJtaej3uuJoIQvEGVXtMyJ/bTn/
uomSyAR6CSoucesodZHV1KkOZq6+Itl5ot49DhD2DQjYVPIApg6z74g584c0kAtni53nkTjgAQDW
4e8lfSIg0+tueJf8HoK8ucztGMwdACujDA71I/w/Jwa6Suxd38043bzaX73NGcumfaRxAugqipI3
rDqPxv/UoUOV7j4Gk/VD9EvuFzwnxgZPlFWcsV5iS9GGry28sfXnswcu51CGMXi7NuKPVUpXb2Bq
YNn1JTke01Qwejpoc7OlOIZcBlGYk7GzZ4GC4OU4nxTn4PMqDk5SMiQYDk9HbCNRc/d3pR3TRnYP
CUF68tU+0gVBf+j65U4cBByanpYVTH1cZsEc6dzsPHSloSvTZvBlg3dU4zzuBPwqT2CKbAMtjIpY
Y0wStCEOp6NianX3mtjNHK3XCL3ri7oP7BHXNlQPcgqS1ohaY9GogA/rvw4NCbHbmvGF5q31o4bc
Ew29FC/EMQww37+6eE20WJWZZRWsBjX82mR6Xk7QQdZ+7GF0f9S1lOuDrukHj3RISLBGEcY7Lc+l
OZswO9w+UzpfgfCs9HGuaFQ0qZWJqBaAqIqt4EW/1XaTsl7qOxIiw+D8fMQ7oq6QL68tL0b2OS/B
WVfQvkTvMFkqAXfJlFotZ1uQMnKKqfr6gA6bVpfcLnWe6ffS/t9jxib1M0KGOeL9QPYSZ7O7gdpX
gBkW8YFsBe77omcFZPVBbxXd8YRAyrqMpMAql7RkHXt54VsSbXRWg6rmkr6NCKG4dlpR0PMNSkk2
i6PdsJ5nFjg2am/jnTCxSBlPhxrVdMpTLq8SkhfF2m3IXwqFAjOANLdXweHKV0O7JM0j6WPJL4fe
vH1sP4mgDz5AXM7/EdHqnuJd5lWdWLrHp+90ODGxVk8INvOp0ICvA+yaFB3Y8n8rCWq1BwR7MjP2
EgZDjXO9S3DNYexWyepLOoqHQfj1b/B7GVWR5e8jSLNQrkBIMlK2wXlqZMIcKVec3gf4YV5wDb+y
HHI1VG/8l+90IV8ZwpX8uCgZw7IDZpK+lsgUd/8LVC2JFbeNtEoOuG7++NIPCjNWYWwGj2Gj6r1h
wPcrqMhyNIbf8PW5WRlqNQVqjfKw4j1khfABN5nsL7wdMV+M3iEaWKtZrW+HcYCQpSNNrYfmq73B
e3XxEEr7RUibkSsmKoJTqA7KsV4L8PqH0idQL64gAx9OxmTRwTRZjlLlsxSVvBc4dFm9CpozN8RS
5LfD1R6LP5FyDrO9COLl03g71RhpKqDZt9annO4IK1PVdDJjztLlTmuFvNHFHwhuw/zkBSxniGTq
7YvbXRXa2iO4Tv/Lr5aXmAxo112lw6+VxogzeBjL/M5KLf2eBqILz5Meic20aV4/L9tWXpI/VORg
yy9eO0PSbfJ5K7bfm9zzPYBOL3q04GMU9sYN31xAKzOOHqmrfndVJpLufiRuN+rSUeQdBDWqz2HQ
nlInOLZ14xs/647I3L6aiETfWEToBeuuJErk+i03WLpUIyx6tKOpGHooDwR3ugHzYPQFacbicodT
fkXECymzk4N6TDFd+cNoh2dKlWtdSEQ0A0Fr/PG6HmT9xoV3fR4XEIO2TtsQ1PRo1/3KFmy3f6Fh
v8TGgXhGqGnL8lV7fwS7Ne+NP2mPeZNAK4drIlculQLNUc+CGhCfM555lnyRKcpZ9Gx8IFGUW8Mg
TNpzHqlNk53zQWbs964nJTKjT4VNnadhECz+cWfRhvwRGbSGZyoOqM/kIdohHNBLJAWAF213UI3X
dMcd2EmoXEWNvehqN9JCd7o0AfoFUx+8sPBMzu3QAf1BOiw+5lgHXo+ViFGt7Jpjg0Mqu7r9SYPT
W4WD5DxaK/mAASmjfCJH5TzVE2UoidrYlHq1KpRfLFAuqV45/mwNq/5YMihAb07IKz/ZJQSnU3nk
EF1KMsidWDl4UUiMmKKlbO6X2DBUsokue4cjVrV1dQ3UGbyrWJONFrqCQVf+oXbOLvuZvzQJ8yZc
wdVn8XO58NwXwvLtmwXZqn9t9nXi/2kuZDFACq6rgZuqR5wpRmOiA9RyoEpC9BdMvVOzUIjPk60y
AiipvYlkudu2HaBSlUZOTfjMTWD+smpdHStmbKFx8lgd2ZFAP4GNiL336QSBI04p+RNAoPTi8WeQ
2sNniNewmoDppBYsHu381aEXeIq75nMspFdyKmwPpiapq4uhSrNhKprBqHNLZPhx7r1dunjxJQ7U
MEvXZRoBd8ApsTf2rHGSKuqinwZtC/+R5o4LzwLNaUYYUOeF9E4oqQx70M4IOymwcWmwKt1/vXMD
UkQNyVJBFHFtrdclphZzvpqBAVW9t8+6UQXp8Aoef5T6aB0/xK3jM5c7/1FqO4e7TiZCYhcyWglT
R+mJEegxAKAmsB7gW37ELTiTUUOtU0sgwaeFmb4S/zT2pb6JShp0T2IpbgEa5WtfCPntM+0RX/jr
bqmAGGPOiBxtCTJCBvtzPPzyuBlWH5TgaD5WURp6jNC50LlJZFT01xf2Njd/bRM0sdYH9Y+diqJs
dUjneuhj4iYqaxwYFAqIEjyDhaKc/FKtKq79CLg6kq8ZA7AePwT6ORXlXX8FLa2jEGt5K/2Zb9Wi
ZEEqJGtdKEWtcDfrybboCnyVXTd2rLNtzlglCeE9tF+OLq/LWvEQUmLie0/LdcQA14X13j4zKs6H
4jspiW0GIuUgM0Yp7jyw9lb+q3Z3noeYeMACWThir/2KpUat6DwABfnxBNRM44i55fJuZyHGzyii
hcQIDEgZAmHZwj9fAgy3qMhMdT5Pub2yXCZw4iVwxWRmlYW4ww9ZD6JrDG4X+qc86VNEPuA03juE
S2+3sC+v4U1STzk4fCYKKsH4UjdpmTHsYumsvM1Gd/XwSJqn9O8shCFiEFqNZCDyWAuWv0zB/ZDb
9VHfniFrSuTyXAZ1Vsu/ABtd/Il0zYrYHxFyss365TX64QXeNsIQ/BVlKjil5ptzxNnUH7kZVkVa
qTWF/6WzXVRS/toRUWvxqJuehIYo7gVNfOb0ie4eakIUM0+f70ug695wIQcgBis/5XwTos0qTUtt
SaETEB0IZ44A/ghuLFg1f3COK2bSYrRT89qkzflHHd205agRgkPmtKPOEHEvdhWxvS1qF2uHa5l9
9/5pHfE6ssAkvP2MixnuHULgcMAjYKXoSv05xvuiS2KE8NGsww6psQ8n+YUl3rEydQrK0nxQFFgs
5JamNijamgexxR1CjZBcV5A5ofGQEAN1y7yW1Qj23/t9CXhqxXIgpQRWvTJIP7G6d9HkgkR5042h
D2q2F239sRM7RU5pQcQ91gIY/vLBce7tZtnARshHODyCA1olcQXfcEDogGxZ2OGMsM/zmNZSlmI8
uxv5KRn9K1IYIiI4UUUQ9ORTerzx7xKZHB6WG13tfDzXYnjsWMLVnPbDEcy9Mq4uq5zcsosoEmFQ
hnKsnLMDFPogcachQDLwosyZNF8qjleLK803ekwQ5Vj556aPK7rILhnLgQWHUmP45moq/spErweY
nixlM/Kop4wmlKgN+WP127hiBFSo6TKtNOTPnzK1ZM0UlxSmWFnUx/olUM7GwU+irf3ucSeCsAx2
yjjTJ/aNLXoeTcUUHufmKhJPeelr4vt4Y1+pQaOyG8mzD4FR4xKLksbV1REWdREAVvzhoH9CVntz
jee5vH3QAS635pckDk+ZwEeqayEgQu/8s2Jt1n1OnqCl8BYYYkdHi7lvXoTx3NNH+yCEH+nqsQ6A
eJcuuRtrger8Oa8MFf5nuGSgNQCQQHLXs+Zhm1xRCOQS9tibuCkVRq9TqZ/1Bw04KtpdCVHYQXVX
cMWPqiRPXp9wRE4cmOsfoNz3xzRyhTl1PVw7GqNrYPOaZQ0Qy0hYy3/wkP0rS8Gw+YcaVGfhBMAg
pvYUjYo6Y30TBQ18QyUQT1xLNpEJz3r2r+MrbVoX23/UmcrKXsZfP1SU1edeF3xfkTXTrsbMTDXt
PkaNmgSy1c5M7IDHQ4IWdeAuVChX/8Kl7sbzkaesDj3UXJzgm2PMQk84/JTkQFMUSvTzt3Ov+gKL
/Xq6IuF4n6V0CibpoK6NOhvaORUv5sXUgU///TxKFAQa29rZNhpGUpJ6ePaiOTmrqSXSynChB2G3
8RE86Q3RhmtBiCRrvU+efcY0A1io5RW+j/BLWSoidScTMPBIJHc1klQzXD68vXC2ayvUkOGluu7Y
vLe0yAP/pjR3+UvapulBBdZKvDEJiei84FvsmaOYcfti53MdCiMNyZbVIo+7F8N/O0+wAC12UpSk
OMvKKQKT4ebXPiOb3q+NKfnXi54kj1W2jKjcJbRIiedaolNli8gSzYVnuBFWUHmK5HM4hYFnLsB3
aocnQYNlgT1iUkinJF0UO5UL3lsDZTSyQ5lmbkU2F6w+vMUcCnZUZkWqQXfy25iwodslZfyDBdzL
Niw3A7c37KP61ESnCj4vT7p7WWruMtlIaCTfC0kDluOHkswbveXaRfPUQaa65pC32NM8wdZnjsT9
kFQGD4Jkg6rD3tnSV/PLYD1eWumF9siHGhvgnopvupCXrBZLbvAfzjkKRsY+4E67/mblWhNQO9gV
p385yCx0d3N+dnGJw9tFAMWjnB4CQEWb0Za7f3GgFs3pniyYykhMPOYYvi9HS7AMJ35p+rCHFzYH
G9Obp1uhMaFp3leMepvMDFRWVqb+QtrDAezej9VWpW3K9K5BEzcaj/IPcRasvWX2R1TehFS/TRBv
wzxI6ZaQ4DuJ3M/xcHCMSf3zV8TUYxOe+k/6xmlQozvqRhe4BhMXDvHtO5wastqnVJVR7ZfS5uEI
VsgFH0g406LrjfnK6V6a4dCpBWJa3aqKCLPpEAg1EiwC+bDNQefJFEquzcNBh2pBekhmyZxy9Wl0
5iJ8g0uOctxMnjjxA4+suJxWgGqO68ltb9mZAf7vSn0yYKBm14O2ny2nHf7CIxg5JtupRp6Rvstg
qFx7sDzAjKqGGnZmQKU5ZcePyzSkpjqfcvIJrIS4ptW+Lkr7iJbrYvbAsuXrj8Ulk4Sychp5fR9k
fi8VxfwB3xisZpfqn0fzTi4d1vye+VuzLutopNZzFzklS5x2x3IRogNuKDPUHhTuSe6wDqwseRHm
wjCxclAz7QecAa8t5CfJbyP3/AJXmOnQZ1iPe2z/29mLLE86eAy3XiXiGVJr0De4Fz8FeY7MFdTC
MK3moyNMQ6eVs+qY0ZkeTBAVctfe0wKBtI1N/sLD7SQQ/EQHZZ8uJ+duu1zY0CHr+34r2+WaMw46
n+b2RWkQH0AyEdJ2cXLWNNFvwdYGW4ZHofDJJni2vpRdisp6qyAQBkW00DH0dw97yG2hkIaJuw48
m2h3AFm91kLLzDEelAgpA71WAEb0b7yXXpBHmBH42XYzrBpT8cUAxdMOkFb6s1mZUe6Ts+LZkVfZ
8WmwloeX/8SsqQ4ZHMaoDouN+IHB2r7aqTgSx6Oi0pjvuRjAeb4kigK4fKimwDyAqZlpygBLRPCe
g5Kv2o1t8auVQ+TAmp6zh8kyFkcgT2iy4fJ8cpEIKy4tpGc2EgJ6CsPBkhnNcHE8GV3T6UHQ31fH
vbwOChKagwoEHIbjlMjTIR65eJXoVHPCa3u5jcBkAurxZKhnkSDs+wfW8UqpvHPFQBKSQ0HYEb2N
jhUT1vXNNdCU2FRaTBXrXlm1Xzkw7HyAUVzzSxK7Uo20cWcby1zIXTnLQ1KrhtKEqT0zVcCzOEtJ
7jyLw1bmJEt+p14Rd3dSgvp+vYQnBeRKpAUNjvcui2wkZLphuJVIr1Cz8FD80RjXI7mABrxxwQo0
mI7qcwcIxPHRlRof/dR48eOtfUldKwwX2Bn358xoyfVDqjAg46p7rZemX2X85A7Tnv+qgkJW9ulC
eBmaRMahSCs9Zt+mboqLtRd2Ed6OvRuMMiEdD1fRB5tq3vzgxwViQ30DtPyl5FLCksrqaBkaLw3Y
zUXq5FRbvwCZNT08ZzYTam7jq1IYTG/4YMTXfY78yKWz1cFskyEYQRCdkCNE3qey4Ss3YeJaVPT1
J9jRrH81hT5gJq96Hhy7mRh1gmN+U7uaRr/WbWvempCHYC7BqkJ/Fyoaj7ecAaSX9zvcsjLVE+tZ
KvKBz93XWeLnXvbJ7RnrhNepPkjGDVLaotTl17GBIkgStWc1RL5eBoGIqWaiDVnLicpf3j7XpMI9
T5phUHwsXZML3YhOqGWg7ehVnTaCg78ECy/MEnXKPpyMr4/9gGTQOMGvwBdtm6hyE7poxh9LLtzm
jsUQoob8UeHf/cgstKwX8mr9oOFoBIMFSLh3CBMYRNvPhodjAK98O2w6QRFZdH0uiBLvfi7V2Q9w
bBsGwk45ubEKximmWnILuIiiYD6DCu9MMAoZkGGTCuwgPVtyIiXEbxA+mXEyL6IKJIBiQaMLmJXb
onWa/Sqr3LwBiq3dV+vmg/DLr7ugKMvtn4BFnEx5IncQKBkdUF09NBpHfM4ce91BUgnkN/XYMwZQ
WIt9qhmAH6DaGB62WV6q5daARFA5sbEa/8vLfMWW1bvQHN/3g8nEj5T6nYUrHDisMaRn033vMfiR
W9P4MHSrADtLp6Ggka7l7W0cNVs33/HuMG1cwYnRMNjBTAUroTPONvBUMD3qQL/rU90jwz1nt73C
3BkZ6WuX1mWeqKxYvX+Q/KvVnXNleBz64dOqnVOilZszAadIUJn6d0b/e30w/oXAID4wJBAXeHwC
W55tsnWh3EbaKCK8V2bJdTN8H1CLSE63XsWlthX+aXsNdk2s/tJBSQAYga0r9rRblfv1XZfgacro
1IV05ZkTQQcQl1CipuQ/HHy4evgCIo6Taswivz/rtAPPVa89SYXlvGRwXEcDeuGNUTdXdThNBFN1
JrP1unNjzf8xQR3BeVHw/OlC1VI4GFQHasrlDTIZALyTZFbo2ZCeqCuSVZhmZ8V6WOPognwwu1tf
q6a44eJ9VquXWIbe0ECQXgdTN557vDN/2JgDoDk2/b5AJFk40lzr1L2eQMQnAK7Sx/TidXmtxCTw
VZft0tNt789tqDg/vcJpJJKLwwGznMjdpGQuaPXz8dvNA31XW7vfRl+Hl3ftreVq3K5kgCTvv6cy
KG4Vp36FrFFOjiMumZclSyVn8qa1h86pydEN02YYHRo3u0pxnjOG1wEPM4QiH1ad6qvgcZ5IvBBW
sRt40HbDtr2/VOSuj3zHUTUSPea2xvLkDISgM0VyISRtZbYQqqc6ytV1ePwYPtE1N6XIkTHlaM+H
Jx9sDQjp2HZ9Vhj1leTJYTpp/WQzbCG4DAOy1NL74E7HMnB5WeD9DMH+f9Y8LiAdxSALsnnmlr/L
R+ODuS9SJF70Yt7JNP/ZDcOFW2dLme/KpMG7QKZBYK/b3YtcrQ38z9FFglGXmhjzXOBGpBzWgiDc
TszRIU9XE3GCmxO04eCkKmo/u5JTga6rhjWSWwpVDdB3zgzhQdFiCahByEk+btE8zzpv4LhJjsdc
ZpYDd7icimiWpMmEyTnUek/BYyCz+2QwMpYYLVKBDL8lha/HB0lu4/RAGJh7ug3/apBtXMOCPXsP
CZ1L0VavccT1ssil1geuoZUiOaHYqWZoqG8mKzBsQuZ95G0U0oa6Wz3KAXV3sPfhrx112TiA1DAk
A+H5mpH4sBXIkOe3gCxVUHBPOPYOU0uPXRoqMIU3aNssLo2qExorlQByrUtteESoxKVqVJYIRUwJ
eXLSyAiNOuNZz3KKIpRnWGxWhefI+9aERDSDFCZ00NDZZE0agRNk4SVbAK1PyRIFOX6dhRcpW8iW
cFrmx7BNda+LmHjzX0/ADd+74IN8+qTekG1nBociYGxgk9+HnKNlokiCpxgOXKaYzooM4pbg7zC8
dOPkGnpzKe3RiDbXq1yURJ8h4IUwQsrp0fZLMIESvfBq910ZCtNYc3d2/JzPMUbRTmBrSYnZUlka
Jepc1yRCN9+gLC9/8x1FkjDGaO3opSOZRDxUqEXScxfAqOQ8vyCQXqmhfbAyoSsq3cX6fT41Pk8F
KgJ1KqArZFUSFvhYihLoQ1bm1FUro0q5fbyExe3ndTj96YIMDWqbs+f5iWfN7TPXjmLEDVgBrp0v
qpW3pFPvpvWJb9V/0ObeGRjZhjvfvboHgwYiFrUJhXrs/9rMBVoUCWFONhy5VwONmxFkKGP4nj18
xkgDF+PszcgucPAi4291aNUCGXlU8vKA9Eg8x4tABkhJMLv+pGi+7IWPDQNPYie9EF7NhRS5WDz2
3aXEkWxVjpz6euZIEBOU/jL20YB7kj7mlkDR+PW5CfjXfKaCdbcQrNTT0V2W80WrG25BZ9/Ye6/G
DfAmKT9/ieDS6ig704nExd+yIJw0Zy5zKQgL4ozCsUmG0PYBz4ZfboGc9L2+VfCE08AmlXljgr8z
81swf19vIszL+45AtPltLpc7IrEmxM4b+DISiJuQFZMWicJJt7QsYepz3HsxKSgCVS3kYbmkbjf6
nqI1bhgqjWeFwkjP4HUFe30AMJXnci5q11dhFPtSCUmxftOmx6+UMNZneUeBwR0vaNLbQZmGvZ4e
kJhWWt7dyZYpaNLCIAxlJJNqK6Z9xkVfO0BkQCMO91lHNVXK+iezK+cal4DL/nq7VRnhnDjdfm1T
ZQxScmTXNhv/uULDiNK8rCX5AVE5ua+EmRJbKj5ISn2Whed6nfpeBpiBTx/oG6yColSktq3k/YvR
tV427g8OOaa9ihWEACWiYOoNUkNeSzCDg8Qp3vO0cLDaC6yAHN7hbTPGxBEXX4M0saLwD1Oqh0tj
n/qB+1l2AGypBQN5N5W13Gl4VjwtkFj21ILpXjaC1lYB6bUswR45U6uI269HACA4FDozwiL98wM/
p8VtVHx7J5HhUYDXJIaVESOdvJo/JoGR5gDTzYaJCnEafOmlkg3Qz6N+JDFk/TWMgMYSgYB6+6gi
TBMSsxa+ZwpTLGimERxcTIYC89SH4M+7lydhgWSU6XYq7MkVNrZvuqmsNxI870kt4D1TYvvMnqlD
czCgn7B5cjqVuXpWBVY9MvkCKI+w3rO9y3TeVOeXjLZlnzg6a5nPIuJE7YKEMkk0PFin7WIKcEgm
/cvEIdd8jqhY3RIjLsfEYMEIRFmnytX9arZ8ZftlPBksqRbCCm/mCzUy05DyWp4KAkVDNfM410Y5
MxtpMKDWBhcGv2YDCcRo61VoE0a8he6lqer0lPgvlTPna/ullnJDvxyangBuVS0pl7kE4GzsLo5D
k8NBUufHtRykvIKTgdL/kfNzvKF4KdMzzXcVMiHL7P0ZpIeotJdRp1NQEsV1MlRnfHlE9UxzwKRa
MDbqUhiIJC3lLlQhmdHZ8UUmPv4gr/CH5qR5DWQxTt83XRvq8XU1IX4CR3rDMCVHk+Zvm1rfLIQN
AGBGGKlH1YDvGQd56Nj7yzTyYVN+hAZr7bfe6JFj/bhjh28IJT1RytsVOAxMT5AGnXpBQpPhN3hl
J8IBHiYddcOpewifRaQq/MiILwm8gQT5Dv0uslFKI67GTZ0xnh3AMWEv1b6dpfsZ51qPKoNDZV5J
rwdLQnVV01l+S466t2KKuJbKbQyS2tyQ9ukzGhj3CDss6E/Oy8mxFtt+7KeZAMuHmOX1NVRnrKH6
Th2Vtx0/kc49pvf8vwVLnDU7Th6oAtKKzNQrrksK8QVckEOh9nQJHHQ1K0HDXqWSVwyphuyG5rEj
QfChzSfepCjTF9uppF536aF3jRxejgYqghyXZZLMg8uFgAjLO4XbeBtSrXk/D2A+2mEW6TRYlITt
KHOg7t+WuLXnRZkyDgknE7KAYtHznAeBstqwaVY1/W+fsXa5MywAaMdsw0S59Wvpg1Qw5TrAwuBM
b9VpenKv1tU+YkS0s0Z3Y9NlJkGbsKCBcgXGndyxl9OhxhpphxCyOYFKFce+SGjQuo1vt+xCPumd
1A2ggfKT6kzJB36nYDxQA8GrzeeR+pmLy29rDfjcuIHnZKjYj3mUoaO3tkRWHTT6wsckxsbdH1qY
gvMMEDfWiqUpD637D8OjXfKpfKvFAAsqZHRfWuHks00OUreXcPAAZFvfSMz1Wv4ceqpxjDTFhZzR
Y03otWf9cJou7sA30l+/iRWRVQZBOa2EtN44zk/DrUunDKuy+MmfoWcIfiQPVUTGnHNJMMxy2+nn
nZaMYyKEU0wqEwx0DMWYPUXf/eDOINp/ybFSJPl1vbaDxNW0os6mjwJNJdLmQI4QU9c0d9BJmORm
t8yBctRBQFDC7+OneecOhYTWIvhwZMnQEjLjo9sn+9nGGerpXEfS6JSvW+C5uaHcFi4KkQbXvmE+
Q2DPvSjcPYfAfNZy784PSYRPzJp98rceVTjkKykk+/4hxIdiBI7pIix6VpXIAn5BKANdiDSByz+t
tann6jLV0PJg0K5fO/SrReqecIkX1CC3B5697vevqvJz8i55WavWwbNKQ4v6AFxiTb9S0VTpUEmd
42uGKAQnc6CGQDJFHm4suCS+Aq98ORiud5b8mVkhBRqe6v5ynk1jTKVdEk+mAGP+b/pLAuQTEWQ9
Tva7Nju0MGXZ1B/Af0cKSLxOQXL7EBPLTWO6au5beGBqMEViM8lFn9G8P5mof36SqemefW4t4f7q
apbWAMh0s0hkOHoVxnXGe+7ue50oyLVSZSbtS9yLUqzlZz8befoB4GG17aRw5VcqlOc1eqdUK/dG
WL2WS7IHgpKT9ZN/ZJ6wK4Q/hsGrxgfzmjRk0r2ULoJdeteDnJyJQfX7Z4JgP8yp3fr6IEcJvhuy
OKiI13O8G47d20ipOXAv7T1drNXDSwJ6qjnNPBMBITt1n+SSLO1HN7/yFYsLXbLDIl5Ok9tPyt/l
xumo9mv/D79OjUzYtdAcJmLJr1ACjKHYLjTiNS7Ibm+Z362ZW4najqFgNun84rACXsGmD11+CpUR
3v2ge8YYimsx5z+7Wk7J1ngwo3Uz+XufaRyt36MZ9WFL61WDAU5Yi3MoVycz5O0mUR80xw0kMRmx
30nGGrURtcBoBUz54hd3p/TDdXY1CfpiCqcFDG7g1dlpOUn5PDmMRDVQeetddOK7yY/lBbxujPAm
PkhMl5ayhqYMY08e3siG3q2/ZF8MWeUuBHWYWBEapSAprvuaVAl9CD2Qa6kmgdOmkfX6KZvuyaRX
qBTFQypDpaXos6Nbuqodvbm2a4Hmg3baWAfIIOvQMiD/bL4gdfxIEVncTp0VgMFkp4tw21nZ7shb
/A6kGh6mVtSc9zsJDMm995iPVlWDGIP7TrXwMwG0ESjPx8YvpAnOdB6VjtYUelyUPayKoSvSsPT6
tp6pxHACuqq4o9lkl7njB8dQsjmc9wjPagZ3m9W9txzLM6aB2RV85hawOl0WzGc+qxw2voZzBdLg
3QdKrBedEK+KSYFO7LRrzHPEBGH1dT6RUxTE4JkTVxhuZhUw7b12+FWqxwxVLrWyVy/vv2UlSBsI
Q8F+N8o8VxErel9SaUFXDr91ESIOnH9JPAzIS6ka6TUGNdTSjJ4riX0Y9m67b51d+OYNPxxrepH2
5MiOmY3G/PD3uh6W0Z8JI2Ml0MojNjW5Y7Uz1bdvHi3hwE4cPE43DsSmTxJ6XNA9GCp7pYLv5BMs
u9i8780Jo04bX//OBOI1lxrHhGaJO1swOI2q/NQDprL84bSd+OqhNK5UmaScFaJwUknRNT086B7J
D51dHp1KfH6tL1l224JZP1N92xpC2GahXpsTgi4kpusS4JRvD0QdYuSKLehrA5P1xH2ufVaMctwn
7iaYacI0YqPG6ZDH8LmmJ/3+GOU/ZT/H/tO93BbLZ9Bk6YDaiLeu0jl23TpnadtaRyebLVuHfBjP
4XI+E5UY6wiBl0tmLN70SungWmer5oj92E6wrC5Qr2SyW6HMVvY74DJmjdrf6Qs8OsF9WavExgIW
ANRP8ZUUhUC/pA7XGyJM7dPvdeWwaiRGWlkoWdR9Bf8rcmZEF5nWXYlZMrUGiVkPzrHxCr/YGrut
vAU4jznu5+p8lKSf/PVVWuJAfDdT6sIHad2je+fTSPCoaw11ufNzLr55hhO/PaUHDvZSWIzSeUOa
liZvVVol9WRPGMRgckVGnZ40HJSgCo2LXvWkmS++Ye2TyqtJ922y2Af3pNDR58z7IIY4KU4JCEsg
VaCBK9CLHNVCvb6BuFvhGxmjXcTFCMDaM1d4YnJ0g21cYAtUM4gW6zuFT6mDTMBH89IQKvdMJ0Qy
nZMbtZ7Am/lK4TxX/SmNjY2eehqw/R4Fsg7eEcIrCrFntXN/4wMYGSSeq1fXbwegjb2vw5SAPVc8
z/Ja3Aq8mgwsqOQsgdnaK6FR4S61o38AcfjxVzWIYEiex2oK8BuWIV0ohfQWfVOgA8fGkq+Exltg
klRQg7XADLrSb8VszUNr2kh14YpQpUC37TFanpQKvtkgkRzUAD9heVbPNaO0K4MzIDpDL+QzuByb
YbUh4dDi4IqqE3bIxBaAKutuEg6IrhV4ArryvMyZsMC9nhD1dTI4ONkkOjaV68bbRUq5LpYmXbB6
Zei6dCO6xpbMqRInUB3FMXwMuUQcH6mckcal/e5LzQtOWcrNxCEH9S+3xUIfHXhWNZmmxD1MXa77
SyTer7AXirfnp3fEyrxN0suovRFY/+EZTdwZMpU3vnK6Gj44Z/tgNvkvI5or2txgeWKePYmLN5Q1
eeXp33HAj9zghC9jy1aVfRpvKhcwRUbL+kmRr6DWdG8vnWicS26GmO6UjWKqZB49veZLjjEIG3G9
i9t+znJdXsUf1vq8GlVxnWy1Ms4CAJSemrosDRFm47jB+hBV3479SVQTY1PAVemwmBv9mC36mEsN
e8Qw5urh8e9bPbqQ9l05h+2tQTmAIhC3z5KRr3qoMPVCNe6fXYGLnr0PK0Ra1YZkYsziq5D6eRlb
kFbPNkDkvEuoP6I/CyP4ktlseW/i7TdZnaKPsgqNg6V435NsVN0GhIACgoI+jxN8lqWAE7l7/HcK
HmIOcWZkw4h/4N5ncnPYaeOoAkscheI2Rf9V+6AZDaDxHa7Si/d8fWhMpC07eqc5O9ZAZHpib1cJ
xMRqIkKq0WjY9jAR4aJUgIu8w2uMvrD3wo6yobhk/+1qcFU7meyZzzGNdtmNcNTeEmExAjl8572z
QIhq7H7TOd3HSxAOPUeJDcei9QHJ1on0LRGckgvrewM+qYwIs9jSnc/d0ReCok2Ufoc1dnh8wxV+
9ORZMC2K7RbUvEb/JgCHixgHWvx3S5sOYE8GuEEP639zmr0Bmi/UCh3aN3KCYG8vHRH6oDJixBI1
6Ulq425a2YPtgk/M9cFFHcy8JMp98Ony1I0gBdoqld5KaAFmWrBOGhY/yC/HydEzP/jbM8RXGL1c
utVycACV+sj19U0isoZQldoY8rYFRvuyGgRkPpVq9dO7LHXJG2Tl4r2uEkLpV3i1aI6VUcxsPrnC
svS0+tffF6Yiw5FsYMRfee4cr4aZRI83m3ivvhxFoO4rYQItC2rHEooR6j6d3+Y6YSzsmcuoA2Of
UXUfLH3JbgT9h+OTP9g/wQWcVb3sYqsJe9yJi2VCmhADeic58PIjtuvZ8GPgIHyHKv3b4zW42GIh
7fXV7yPvjGZRn6w3HxjZ6Z4aaxOWPoHvFDahvvHZWpk2uXffa32bH7c5sxhjNYqpXoHNSnp85z0n
JzQ074r3hLcjVKHKi6Mjd8rWI/F2qhFyvEKlq8lY5izRqP3EBPTtYlG20eAO+AFnz3aMyEbqt2Cg
aXoZ7CrozPoNmMHy/1zEbywiAcFj9V92zVx2cXfBhg2RSqx85rpK/A1oYvZ33XcOiS75mipjdSck
XJ1ZEHHPPKskeHjJ7/28QzQVb/Pwsg3Wvoe+ElhsAlumP9bNH0qbgqz2GYfz0ILAsIuqgb7Kc7iz
3bY6/lX8qr4SZdYnsv/EKfIyfDEa6j8dr4kxpKZt6QlaB5eAUvlXNPib0x9GRMWiMrl5NHQTXJkm
Ry6kmG3x2zAKPzxxM5KXND932js4nziAD6s6b7x7K0wfsVGiY9GKAVFV3unCp2Dptg8sxhQVbLKG
mwNU8g1Ecer+IQvNTB+ao4IskYOSKaRHHLMEyrsAek7PBR+HpqYUjjD0gHmDw3w9rUNtT79pnQmi
FoHDsYV9ucbZrauGaa0SIeF6q9HZxDT939g2Uw2RV3yFcENKZWWGkAtWhm9rWEua9e0zitX651yd
+3TeHnxTgz8fOXyRTl6nNK+4lDUIM0S1MIoCpzlq7lt6NDYgyPp0oZfRVROyUla+1O96DABA2exR
B4oJoyJh0J0LDqGukYrxN7NwF9RvWnzTsOA0rygVhnyR8U4ifRqQNrGL4Bz+FofgfIJ7Y3J0jeNI
sISa+smzFJn1LIrjUzMnBFpsjRGXjrD5qN/6hrV5gaFxowjZAdQ3v/RAVi6v1AD1TFi+5giBVc5O
maahC4bq7YXVsxfUP+IJCMsCopa3Pn/80Bhaoph3pzWtzw68pVsR8jqUDb2hXw5xJnHmNLLSVMo0
Vzm63d1Hw64coFcReUHQTr2Z/obeDT9KpB9i1BBNmOhRuGqGH5iP53GMFMs4Hmm2AqRctQJE4Lah
E01LXk7BDwsr/LECpgPRQBwebNNNgkHPwMDEO21rjXSL3VnUWtGr0piknGC5Edk/Y8l1YDqFIfRc
W+zJazCpY9M6XwMjBjmdU6c2YfP3lpBzZPcK7bMmvYFshtcitM+319BnFJeRoZav8UiseCislRF+
J1Lh0aB/zyofMOsukL+bxDoMer97WM6TW83Ka/K397AkanG1Xn81mtFK3ETrSLXFzvZBduE7sWlK
kt806V6GDkXgA23T3zkJI0liSFHK1IL8ABhrw4SwZl8hv3mH0uCK1oL13HaOLMtBlb5vjKS/r4WB
Xuo70pgpKCjDgTnbTnjnMsDVtA//XVbPFKwg9q6/4soPikkuFcW3mQfLtLXjCPbz2AssuFp+mNM3
Z1BXVOrK+xM6re/YsMprqJuXuMZAIDtY6w/gP438EGGNCrfPeA3AL5e4JFIlIuivxjZUnUOT9UTR
esBjss4IsLLqWoR/EimuTiSU0X/6zANxOSxGZnNODElL12vDhDulkDVEIIccGyVl2hJBLwF61g1k
6LYswuhlIeYG6aKNcbqJcdwU59S2zsypgYXsX/nXwJ8h0ve+MzSb+Kwep0ghSNQ2omYyu5J/fHfS
vka8WK87AzAQZmXyGFrrhntRIUpsOAvpDamOsJ7UJsG3MnyPJJEL3u6oX1iQzooXa0r0LzLCFeSI
cHxK+HB9QrxtASVL6bVCN3eH28Mm0KREaJS7lDJWM9cTAFXyT8+JewwYGnHwqp4GvmEdg0aq7iS9
30nf36B0CrhoR0SvxEfBDrdyTAFPsTzuh5rtE8kaR4DNlpCxvxIczNudw7rViacgvt3k/G1xdsJc
tk4AvjYmJpys4VjUC3MNIH2O9Ge99KuYTJBNGfDG8LzzJTLt12+h2XzPDjSUA2OKTtiCivsDj71k
T6F9Eb/n77ksOLeqJrULKZ+Jwag76Bdul4/U62gFChfF83ZKa2PAxMLVDW54QkdKZeJj+hcD4bXo
lKUCyKI46HDpcmpx5BxpsINfoVLpbD48gteB4hiNvExRPxAIXsLGWqPef1fzllsmjBk/0bgcUpyx
oyqOg+D0142Zc3xzgqkaSk+4wVSjhbwCEIQOCJPr5Dn/p0/87FtISdaM4axw7CE1qBvyg7u/0noU
XaIOAMsrGNDtQ6tfGo/46n2V1zezE27eDbIx0zh1HE7FHUggHI89Mje2i2B6NA9QyqijEu+KKepF
CKtmh5W3sufw7XsXG59aZlV/EM/7quaMUO+D2/sM+Mc4T5mA94n/+GWku2/dAQS+HIdCUlLXjmDD
4jec+ryw/cKkvzl85SYUxwMNXO9NCb7cv9M2PhhUCkIneyN7/11OwwoOgDAX5/XLr9qtDBWUpg9K
kEi+3BBtHO6yxh0/4Tqr0WcH0TBzftXxcCTQtszzSRhqpEVEHQ7rOupc5f/+uD5Qtn30LfN57JRm
T4k1aSpQrDrBRG8XGTBXfrw67ynfCC9ee//0tlkEUXq0ZnO6EnwrB6o+RQPiHNSAVC70ycUyfk67
zDdwc3ru6OK5W8dA0F9amQSe5yGpdEYpqf/REfTKgKZSf6YfUuaZXj/Mw8rKCe7iymFEVKEuYaDi
URu6FFf0oAZ4HiXKtmpdReP7AsASeTLjyD8cmUKX9tAqS+3UilK3M0UDaigJB79QDKN6Ogq8JkUd
TCouz5Bm7/mZCo8qpjGXK6q/aeo/bBnR/zyTdivh8FjS7F0IlMUPlSKoFAZATOz7vHL+wM5HsZ07
8Nu+MBPD6mTtlGUEAL/E3aoseRe+9gxS9tMaZ7c+ATdP3mI23TtxkzoZhcM74/kLOHVBaoBAEQRx
zZcIfKGSt/QNboKDCmjNVU0lLNe9h60pg1w6R/jM/lqc6QVRomj8zTWf6v5HXCWqQICWPUvKhj9P
aIaruGXUzuCukcVt+9dYJUoTRYT/25cLK0TDUwQwe5bR3CcJrF1U8cDp682ikkoAs7tcVTM7ClFj
zHcjkXumT2e6yY2hdqwnhgulZt6ZGx2+rK8mucdk0Fdwo30sAlnc+jOqYJDpIT0DBIaglXOpfO5L
eN5ziPjZkStlkuv2m9QuWFw3nk9YnmJ0NpQvt/mCJjlUQuhl2EUvSssRWvUitqq5VsOE+W4H9bvU
hssOTXZb6FcUZZoOqQhfaOf/0LHTsgwu5kAy7JDGQSoZtPCoBEgsdpSDGLpu+7Z6sr0y7s4U0GCE
5D8Dutty9hNb2Cf7xmFA9thZhHFwdO+JyGGP7eRk5ZwvDiXr1cxLnS5oG0Vnh/uPioxe9kezu4//
/6tQnw7a7mhALJgnAE35g3STguip51+SaILdA58QvWvNqwsB31onVEX08PSNIzWu8NGeiBNdM8hx
vo6RZB9N8weOEkdZXn2Ia7fVAH1k9Xtm09i267wdY44bw0erZ8kgjdYKrmJBkBOX3Nv3U/LsgSR/
tL1cxfZ+A/zb1GyIySMo0CqaDbUYCb2jdMrWSLwaC9tkqNp3g4EkdPqPZ2i2gl2zSx91vWpozKwx
cuXpq/A9iYr3UvvYx8B0xTElcKKSb02ebEMTu0/yALLEFKGaUJW/1wZYI/fAtnxdFNiWyL6VmCAn
uAvSvWrqi3/+Rtj2OgYMaCQzsK0FCxLymtzxx/PQBA+wazuF7GZStl8QiV+XXtZW2guAYDyML994
oO7cxupqBBAx9inByUdzj08xFXMPU/GxVwNVhfOoAQ9Dm/Jzefrq/iloa9qKzuusnkMGaqo1SXci
jGcp5pzucq8iPV7x8d63rUiFVAbCd7vPXgrfUJOAW7vAQr0n0ftg2KTHIivDVfkLuLV91D4Ds8qr
5g861SiEhm8BuIkPeUmgBMjXwAtToyY4JN7idPsG+5e9qUXZNtKW6rHklUj1WL1GohOZMAU9lpdI
DDGFhjrUH2u7bWQQwmvR8SOF9eJLNUXH4nlXQQtPH13/xUpmOhLq6ElpGmfn7hF8MgjGg91XoaJo
urvY2cK9N/Nye1VUKnVQtOQFUiDG/5gvYaYXkiB/lycpr+UPc9pMdm7XbPabLi3E2cw42ukOxEyf
mkKu4TMVsjcexy4g2PG1Dlcac80jWLgWcfCTyGptXOQFAB1D0xgRSmNyEKJlu0k9tG9LhUwvOrkW
rvy3jWJLc8DWQQpbB4/AeMmGxDQy6XArpRbvsY0R7Ur235uSbkAS687LGIy0vGK7n1Axyw3HxEnC
MPOPbWyUONh+ytEZQAQ60RWXGCkedzTLE6lrZmVezwx7DfdzdCdmDVVS5JQUeczlMeoCcoo+AoUY
XStCeLoorO1IdmAX3n0Clsz64J7LfTtcKQsAZtUPrRVnLBNQLxGjpWgyLfHOYb5nACs9epOx+Wj/
mlcEwebr7vzybrgU6xOBSjow/ZJ6Ht2XmFLB1kYmsYGvHfjWW9kEqDlzFN0o8yl85Ed1+o5Uwj8z
KJnND1O3LyeHlLBiXzV29MmXmnkgyjLqmKfo3tH5na05tS/lVfdwZ8ycLHWcnAJBgcfNYi5h0rFm
E4epzV2zAZB4V8sjytR+g6djUVTRLs/1Q7GTBwRXstdBEMo65VKQ9THFxhiS3EKDt7Iw3pRTlaDl
xSx4SzTe12grp0sRuC0KJYAOyYLTFRnSNdnUZ4uj97jINt56Hg3SmI8s1eTTu3xkqyZSDqVDrb1f
ghMRuuZ9NoGQC8lWP8otrBaj3bBYO3Fn/OEQ7sWp4mOxPu7H6xBB9GPT1lwL+SevoNGOEC6JzXTf
MJ7hsmxDvSxCuZi+pV8AQlUmWiwBzFZ7w5tORbxTZZseXE+h+MkpYkvJhx8MEiIkgGP6XHLIjB0n
4CDDGL/F4qcxpA47q1x3vrEoxxVtmU88RIrfYhBjQQK58ur1IDhm9iHUeD5PXuEHmlX3+6m8IXrv
2PWQG7Q0iJHh7PIhrV0TEYxTCHygkW1DuIFCF1fWI+qBjyh5aC27YoXI8LnFXrBa32mlvbmIeMpE
EM8eazS2v2G/1SY/Taj6yINcW35uTvoV5aj+eSQ0srL2nrx/8mWSp6OYTaHIvidXBKmoB9tL+e5c
Npw/Unw2z7CUrMy+pC0gLxK3nsCg6zh/uN1RtaarLTtCRyxg6T1NArElUa6OXv5w5PUgFsgZcvP8
u1mjmsNK7X8k624Iq7XAjrJDkV43lFDzR6TbuP9U3hSdtvS1ThGN02mcYJlbNjHWfkRFtKmdWKAc
nhxCliukNNtjN3Ijcb1Hc1BbVs5Ihk7P7vpa0hH1NmfY+5C+idQX91WnkmY5LHFuYdyW6i6bJnOq
WaARWVU/NY6IGAPq7dKKD1Q1VoEMDbdU7svy92QRwqFlPU0sXZVhQbhtZ04iLkvwH2MPesyo9qdn
2gzRp1vRxxwI/ha616Fd157MYzRP1GZm4MTurE2FVY/NcOrPA0Gw6EN8wpnND6DHhztZf6L36OY7
8oEUN3IwEuJhkPWHR2mzhB/THwX2rq38J+tfuIJuh0yyL6XQwGPDRh84F8XqBa3n63AsOuqsfjkD
VYLMoUyXRwIJtGnhQZxU4ccIYnHohfBoD3W1P1fMNCWhYjYlWpRl6a7SspXRm0uKSIPuZcxpEADH
BkUFRigVHmTQXo8ySIYevAgv8LrNu6+IizK23W6SWE8LtzJjdeZfZCp95pNBE4Oyf6ymkekNavvF
W+5g9nuGBEATGvRqskA6w54UFkVxWnWPYM9BeHtp8SxTKszibvHjH4lbpevynKIUFAI2y4Hl9EFf
BvJUTnDEhz+Ppxm/Fvu7vVjnIh/syviys0A+WxfwD2vcPszGBWBuDK44NpM9TRDKrwZnZOjlQp+T
xH/xTGNQM7mzVGuA/b1nZR2yDBv64RJZkDQTehjW4chBHkgazwvwOpXCjOlxu32xVF36YITir9p9
/FwGTfBOvUhU+YEuZm4UlZEJgGKSYG/khc0JS5x0sv5DuJw8Tz4rEKJzEyS6oip2eSL+fZhOjAfi
19drCjjY0pSKZbAYFkKBp3wHiCrQfz9PUV7qhV8kWlh0i+QtCb5ULXxTQokZYeAZcpYyxwjYwuxi
zt4Rj88TQMUSFl8TQhK4qVqVMfgNwrrHAKPbyMdvJx96rC41o0/jQitwYOK1NTOBCem7qR3n9pVS
cy8T520s1Z/1i/MYSsW3U1PnSW3P6DlwzEilHg3Q5m4oy3gj4M82bKEyGNU26149wcduvwCX3vKF
0yw3kmdetgTkg992FogaojOGzBUkSAfhXJ5wNzrM1sFXdujYCh9c5TEqrRiUBrAR3rXRHUYI+sXa
AOJZh0GochbGDA5phGaXGT3niBWPIpUux16T/q0SiCdGjgNqNBD2Tt3rZyWCvFqoRnby2AVRpCd7
Ul30jAwjCu4Zaqys5ZiOhFRpUmsEqlsb28P1dUPFVkX/qCUOWOa12JYYz08WJUkSO40r5G/LbDoF
bmJOUCWL/mFEseg6d8CTb7SgJTM329yvGdpaZ/2vQ2+LSu6m1FG/Gy/9Xc6vu8/VFXmoEJeRAJrZ
xvf0qSExnYunN5c5xu14jDPW5/V057DxOISUOjZbe0oIO/pEujohcVg4iIzsCvqMkH9sc8gAigX2
8OhyhL04tOsLX31Hopm0QOWBnvg+kYqUlNGPcEsqNx2KxIWz8ZJhuuD6NjWle1cgG+g12wjYU0e+
rjdpXhkADie9+Zk8AS+ijy4K14iuHxMcWGuNBu5PiK/IJaRUCjaVzNEClOS3JCi/XCAaJJYqozk0
dRshEeHFGjqL0SHu9/vF3tSvX/F7CF9tCYvKhISH3POZrGBxIjZfWaig2urdb5gNwdr0wQ4nFd+J
0cDixpiacCqISqD6UJhH8q5oBNXapJwI6/PBpKUvLY/VSlUZ3C+EV9a4KYLNIVp2bfmGFBgp+kK/
YmW0yszvT6EGx7gxagtsSeFJvktRWSJr540HDzTv1Zf1WHznqxfdA9p0ezMdP3NCNRPFeLsmplaO
abIqbd2w9JCjuCdjvhpeOeat/CAum3T5Gl8uB+O+fg1NCPEMKitb+LJkRCtTt29sbhtXH3PUi2VU
tj/6qHuhjZTqDZp0iFoHyLiwlzD3cX1Mhd0dnxxm03EWtW0KD0fg5ApJqO72Vz7GkuZ473X3iLMv
PRm24RijhfWxtLOk2pp7T8tnYTa/9wUO/wBWJf/AcfZ+zbuSpOw2v/ast4lmIL/f2y6d30AYZ8qk
4LVKU1cMZvFJP500DY0jcpixb+pAz03lN+9Gc+2WeHmUjEKp5J82RGoa0STxcQFT4/gGWG3y4fgz
thvOzrNZoeSV1ItnK+gXjgw7eapsyTRONE0UvjfnmGg7F2nmUzTHQWXbKMQs0xs84/c2wECwsYt7
Cvgn4kwepnKhTexVt/wM73fedRMEuP+SfsJqQsuiky6DeRwNRhTb/EBu88jvPPfdR3r3AxuHQEmy
Gh6rFnQe3bDbaPpHdb7umG5PBMGCegZVT+EGMH26+od2m2tmiy/A2Hg708/QAa6gSK5kWcSmkmyE
Aj8hoF2jbX7qFiMYE4FMY5rQWV9Vc5BMzcIaiSKjmDOi1xTC1iWJhtS1bgsoZ8KNPfvTzZESmMd0
rw91mut65XeCazFZKfOVG/b9K2INNNUefq0lpt+XcE/q8xzidKGQfN/UvBduLTYB7sPxNP9djrtl
pXPzf0NkR0G2fjp2CQhtu2d7Yw7orxOcq4qHG/n3yqUxxBv6cWsqHsCr0r82/1dsMY8cOpSFBd12
mbSxiacq9CSmQ1TNXiW5CqhjqobMOSiIBc0yn6Ea5u8OnWz9anPsglntn1+8Qhj24jPvCfteDPw0
ytgVhkMdWixRbJ4wnGl3dl++ii8TmDXEK+IgTHhYj/RFGHKxcaDM0cTpzcMh91t+1AgTCuIWSz6J
bJdMbd7aNjqOY25ERPXN9FZtzfu5Pb/trkqHSPIhl+Kt7x7RDAxHQN+fz5o8mK5owiT9HXIpY7fm
L16mIaMkCUQwGOccK6lwLUTZTkI0nLny6PEHdOHMuD/LXYhq9+BT6eR3YmOPokMD5ppOA4eFsZhw
0HrZQu+XSQDMmMvnrkRGjnytszC1MdlUJ+zfrvwBQvfDAEwtx+iNUPMDYQBjO2y8LxGR+DGH/bf6
ftxMP6qbjTqyiiQlJrz/C024CtgecpdTebjjtOm44vz+bOdMpW21Lhd3J1vsjt9awFTwi7LIZCaZ
IRLLXbiHvhmjL1aOwtvEmbYovEF5MGG0jGvSzjmVtwWwTm9/jXmt99hOxVz4Qm4MTK3xuFwIeVbn
lqOrIk5q5XPneb3SgQ4151qotPwK4jPf7KxLwVIuAVzX1Obcy96M2cxGzE9vUFF6TrED2xBVxyfB
jqea+D56er/DG7iRp6QFdFOxylMANgxrowWBMrxX+A8FschYcDTHKDYijRUuqtDbPgvUoIg+09No
lkLKSugNCgMAnuS3elcsXbCUZ/w/niZuYvsvCDjv0EBEbxSES+CfW3d0+34N7UZJgdaHJQdSXKwF
zR1r74l7lNOVZlOmJUvksAs+8MMoseYO2Dw7090Uy8DtlNuuUOTd/6Pk7MUfbW+VOAq2i7rnmr9d
BDyVg6XQ1Z6OUUZA/eUV/jnQ8QO67dp0q6KQnZLIrWBvqP2Ar1IhzZkBERln4HzJrha07hcP+Atr
oTgAaq19uaO+uHrwcLRU4CRqnpCv+2bmzD3tJ4dUBfLz1LTqSD8xM8dMhZ75lsWnwEiI5fZsg277
zw2buOl8Qyx63yZ1q0jzpc37WOsB6xM9FSi1Jx8mWfl/i+U5QUa86chi9XjmRBSezJg82DYkA0w7
4m1PmsOdT86ugPIyTmOz5dFB42YVc7b87aCkQi33Ab/yesZDs8bQFkONivvJtspTMAW8741kSTSr
TnyvdP+0Wk8ZoGUkoe3YA1l4XJIE43z1yKSR2r6s7V0mfP9u7Mct2CBzudsVgl5mMr3J2EGVphPA
yVc4oPPoXKsmipYg4HOjnlW4htkKUStSGg2FpaoIb+bpoCKGUto0SmYP2IpVGTkBYXi6J98tgo+K
G0AXEEH6s7O4rJauY+3nHm8984qk9QvR/Of9TWR8ia21WVKRIGQdgnSHk+V1/p1UpzFm9R2TsxmW
Q9OPHhGHIEdUKIVFcPMb6JRY5Wx1VzA9CfmTEXbbB22Zq0ngLPqz1TAtS3aqxgCiXRMZD94i6Huf
c5w9ME8iXSGwbDo4cu3ThJ+qy11ReZOkmAiY8TQkQ8uQ6Y2sodrPhWYRA5nYL6zY0RcNaRqLAf2v
Iqc2NkjdssHJL2e9SICp0++a07q9cFLM9o1Ch9waQKl3/BRQ4/H6d0oC/HUaO5ma1hW+r/Jlh3pE
vnb7podl849kJ5cxGsFZgVV5lBU/2FDummUdH9Lt08W8Du3jT+YG5QlWKB1exIhHR8jAxUKwoXjt
y+rpLkRAckxMk2JeuhsbWtuIziQIxomeLTbayMKyYufs0oVMlV2IgmWjsRq+8scF9BwG7nBzwwcG
1ytJSopt1GsYaTsg50GvvSz2hKVhZgoqGciwbKvudH6TUdr2oEnNktfwC3+ryIZM18A6OYxcsDiO
6aojSC/wm2l5dno/vMCTIwb9H2M2cWyADdW6YJIx6jJwyK07FCZZSSmo+5j3KJZHMLwTDTBlSNwE
+YG503GlASqRXOkecCXbOaSlT41rKkdUinlaSsv1Z0whwbVlfT58UovGefwonrNiaEYgfljVdBgF
xyZp6+r/E+RG13+LcSU1lBQ3As3u2ZnoVEu+bdJENwA7pg52AGr7oBOweNY+VRr6Fsaorkp3pv9l
2qP+Xx+ldibLUfAlBMRIw9XHgemF0Z1JXhdWG7hpPTyELWYDFHEOc7lYPWpfn+SgxL9WkYlTESoZ
SKOgVQe6Vy8Eq8ratrwPMdUfLyi3lQDtGxfxIksGx6NE0UcNf+MYfRzPQ7pVl1yfwtqzFrRFmlDk
d1O3dz3QkqDXt4KhmPsTuYCvyHB/bj/BVZqsucnqOzENRWta4VQno1C6PQc5kafYk1HBkZR6oiDT
FtkqXj0RUDAr30e+I/38y6nPupL0C186DiFpvcW6OrZrX9uPL8HrLjl3AmnRv7SQK5oHZYsz4GZO
7BJOFc3qnu4l6GjUkef0KPhRKmuoObd0j9UsS2VHiG8eM4ikecHc9PafinaQQOpcuCvJz6Jz38LJ
7b5sxv32PH+QUTjspriIRL8mFApZPZvJQC3A5rrlw1SI6//l+qt7N9kFf9QgrF32ssqvG/tKhcmR
Jmwju9mgUb5wELhjAPmoGcR6GrKUUhDq5LDm56eI8ineU47MVi69/uJusx7+dM7+oFMsEPifM79g
vW68bLGO39o8isiGLuFu/csADe6P+/ZyVYqKvZR7KGFsDsxY0+VRgMUkojvCD5YjU7B3Q6+O4hTC
HNd/N7LwVoHw+zxts5Dw2+NYFglyCSV75HoBjx/30rui9eyNT86J02yPeKWm68PTi1UdXzxhvBC3
bCrS+gYMWOEOK9LfbHhdWWU4uqz5sbgL9xah3qSBFNIgxb22WWHkeGIX8X7KpFOyTIvrJhlK1Jog
UCjAihBwnvIhuirP42OJ01YeHCZ54/mbJLo6GIsDXt/VwiaEvkxDFQ+hp2HuADVmCISpzw/XsRon
otogqKXJUyc32e922rbn+umHx3Zt7hQEgn06I4cOjlXWbupUgIL3Rbc+dM45aeXanFRqIk/ohRxD
6O8owSt3edYDJk7engzhiqS5PLn7N1TKs6PU+iuZQshjP4FZKi4Us7Ryl3GifkKwqMDc36tbzyUi
mDprDbe08akAbL6ckR/klAj6g/cRigJQ0oujw3XRhVOwHLWpqSv7JOA0m1yHDCVI9cfNhjxD6qJH
jb3fZ8QC700hvsCVY9FHwEbj//WxES3tXF/LfJO4r25JZI2eeFio8dsWEiAdrT+reJswo8riGWzv
42EQ3QqitbmACfLinuJdPgxSfqR/qvDmwmjmOimUCTZqdtNfAIX/pVF8aWt/j05AyKnGiLoNSAue
KpTRWGwqx+buzXMveQysLvhIOzTrv0fsWr/XdpsR+dtlGknw3TT4cfqxCXEg6ni5NU6w2fZmFD6t
r12S0yhXAqf/jxC0hAuxbpJha+LTDN+dm01531Kpfn1MC53cEUyOiX0mI9Sa5kMM8pFLApJOKdeM
dFl2JrzsN3fV+zqu9hmcNPXlff4Nv6Q9h596YRpgSVSoh6H124M2jMPJv903LUKlDeVHrqGuoFYd
sJzi7fh+ocwPvYedP9E2gPi+uhLj5NBH4XOhVd7s7I6yIm01YPiG3BbmdfQ+T6qUQvL1+ph8Eyyn
mrdlUY+8kPhtSIuSHgd+fd5osQHFlECWihipCnyZeiBd/ySC6UGW17croFwKZRrtJdFdR1wVxLfM
AgHYeuovNAeIgmabVlPIlvUkGMfaApM8TPZNIYv7rKXPkBWxtD89n5NGc8qlalr+QlwWbELGXehC
cQXGjVF/pZIlvtyLgwpvfiYekXWUk3f7qGeNGGfNpKog1xCC5FLkQ1/oypyLVbspVHjbjW3sLL8J
XGJsQNGjq2nt4ZcAwD7LGfnX+MSYEqdX2Aas6PuBva+oC/Z8xsLB1EF50Ge/s1zB05Z65IsUYV5f
ZaCRYb0rj7fNu05moyMS3CUeS2sQyxHMKnBsIRZ9YNziRydrnfxgiOVn0ROUq1d/CNRbLPyJahW7
8vk6NLnm7C0q12QYAFXPOv3kdxMquKdvyOOstlfLcPRPE6n8HyZ6k0Q1omrHFgGMr5C2jxOMO3DV
bXp9LNqDfIAp2c+E6DhX8TZokuWHKRLDVmANL6GzrnvQNLZD4Z8xHkn8zkZuQL3A5p9jErYeFSwT
4qmXKMeOksgbcObroBtXJIWNhWGq6OQvm9KVM1s18gIicUhhErBw/sOkRBjcyp+vjP2xQd5RRXSC
bK0eFnhNJzD7onlwPZeSce8vlLyJ9MlSoNIYN5XhLw3f2kFRU1uWtK9iuSIT4jZo1SLnHveSupRT
d4cD7HmFQdnMPsiCSxJNBMWEFJBzIOLyEtzU59hdLtUQiLQpPo6mBF0DTAyhAf9fWtqpZ78JrqjT
5dHGN8WBL1gRUP4cYk/azzEaYj2pq+wcB1i6bV52kScW7AiE3pNZl3V0U69gTxH1DTlCMTGhVsDK
We4JrQaOiJ8Zettbp6uqA5E9ip6mMiWOJLPX1LN8hkOezpV5k04HfkdxoF7FoepfuSbQxUmF69D7
uWGR7UB8woA/r4QDLhOPjrF8o6LOCAJVDJqu8hdX6AHMqvSKHzvk0I89T5/C+k+dBM87BVJQkkCE
VMrLStVKq/MGa7Zor/+xStH9uC+0prKOvSgkwF7OojwxX7jjG6ZSF7IyEVO4+QEUEN2baBZLgXCv
POkXZhYL/zylwgD45uI1JMQ7vKhWEScEFHN0vR7LTEKNoFzQwFkSFXP6fiAceWnxCsvt85SP7Fe6
qrN733W7moag/FUbstGr3jc6Sc4bGBbGcSj5DUtk7OYVF8DImtUfg7tKzauTUTId9l+jbvZFCVb4
iTLBDiIIh7/evc+z7J7lgyYOsm3EJ2qAzx0V1MdI0BQ9D7isUrQFMgd7bwUVqh/Yr2g8+QDy8zTZ
tLu3lWxirZ99Msk5J/HquARBpnPSU4r1i6/h2osUGEWjvKc9SI3uIbm8Ml3wEbBHTQkHn1Pv1mIT
rpm8qRstMuOPWjXRUIywxbDuL6vKXCgVF+ZP9vq4UigGiGqKIfByQrxBZrxlkdEqNFojPTh+/QL/
kqBYM2oks0Lyy+V123RqenFAre8TjE7LuFoVJderBgJs7t/Z3C357CNj6LRlAtuZAZlGgf7iCwXM
Mik/bEQJcCpbLHva+JmxCzqzPLpK6ISmO+sTa/T5eJIHUW/h1xAGHAEoqPga5SwFHa+BMA9cx/u1
WaWuhrBR8eGk7RNEoAey5+7DM3Bk2raKVwITr3eUGRfdinkU6tgX9uOOwKrWtBdpaanRK2Sfxdw6
pRXsvM7dC5bfgnFTiy4ueJ6rjO/d+C3uFR0sRRcpTqSk6SFdolHu2k50FUmOSJ2HrJZL13wK7MAi
sqHyMXLUHqd8XH/h6gIW4TiSqWpXYatp7f7qVRhC3MsDM2n86maxSyats773OsZ9n5L/1oRMJyjU
9ugu8bST8g88Iy4+a+BenuvqeSk5IvQvAlTgisZOJPvSnVLcNorJXq7DqEaWWlIB7wkkE3ws4/+y
GdktPdX/3cYiXBZvzty74ILcATgNBZePIK7IXdhRjRA3D2jC4qkaTnqyR3zvJEstE+KAhXKqN6fD
pUMtrwWR24GUmx1m25cfBY3b3KcBatcPx7VE4tualatSsv3pmqCgWnsLpChPpESH0rZLLeicPnH+
9SHrAln5Q1AbQtu6b5a7cgm/qahqMfEzB8HSUA6WVcJcb779pkmZKj2U7Vbj3Ru4C+ZMAL0f+EMQ
T7LePt8GJa9SO1D57Qhw35ilgL5pUsjgF0yNGTUnkxqwJjy44hjgsgGrYnE80ap/WKVeWGfENn/i
8yLxWUYceQ/qnRRN9ai5rMgQZu6ivj4yasoNGxN+yQZa61246Lpl1A+vAqCFtCeFCso56OnrYnlT
QbiRW7GstIE95L04+3gO7ePQQIBS7aGY89aoFE9w15kU7OJiR7VwNXifAQWV6jGOo/QTeEERVHUH
fnQ5VIrCXYFg8Daa/MVY+v5BOM7vyVf44lb7mCN2yTYfOnKS3VUMwZmuFZjy/w6VQsTbKmssI/Sp
zoFVLMJto7PXsuPfuAruqFrJkmMfAkNxJnIi4JIoE7Y3yRIGH27CU+f411KVzHed5JwFApS+B9nA
HYv3Q9h09sBnQX8BrmzgZ7dq6/rZ9BX1ODP32JAkspyOnFrV0sPOdgOVbripfUNBupgzj7B75poS
wmD6d4EwdhGSwcUZMDVLrvbfhQsNLimVrwod99KhraGsG6DW610qfDA7JrBJWdFpld4ngcyvO5pH
urpnsgwi2cxHrAlZWSkkbKRharM4/Nnq/qH7KyvnZdRG2nvUhNbllrIbibU3onX8JO2YXJ+q6CDq
dW4nGzYuTxVgryhlvGU1oGg7WdX++vawfUhdvMS8mrZp2/dKxbfYY1XcQT/WGRz0fzhfzRAK/oMq
iSeNw2PXKyowrso05D7qwd21CSb8yBPoQ0+ZuYfqvo+Y/BR15CZ5xLlRWkQJ+qrCEMGOEccbaEtH
BuF52CvSVJVBmqPYeThxdjEry1iTA8RUpgbBpaPUg6UdWTrQVQPbKgoS79ivaQj7ra/4yiTSEVre
o6ZHcQuQrQS4eyDyEiqAj7J25zNvLc1lbYrd59NdBCrt3SvFTYjLr8DA73ejygQnGlgGr3pe17i2
IYq0ilFfhhjjfHsPtyzRObRoH8D8Nj9EDUzbf/K1mlJTVXHQy8gBoXmFlBDb7rOTVgKEqRZZ3knz
UEdUm9htUQRKXbkl6T5eghbE6c3OALhT7NjTNE9CwLsfFUPC9UBqFWLaahGs6HURKoxg+58NF6SY
iKSbRDGZUm/p5gKZPx+K1x4WrwiF/kN8BR/oqW8lvVxAOWak2Gitb3y/uKvuUzKdnaiUBok1x07f
0ERQuEp57j8SjSXrCiZjipVLTJ6R6x3APzoCJXMT2mYu7qP3g85Zm5MBpo1nRA26hhvnpf45Auk5
326VSohJfg8II7AMiZvxit3ed+fAFsMkqWxqz8Cw/E1yD9z8Wub2Tkv+umEmDZF96o34zBdLlseL
mpXaHM5IpOUnq1YYAkIJfEOnR3cpbGRamS3Nq8ZWVVTZsXfuInBz1RFlHC2i83yZjKO+LIhcyNBe
7udXZiaMM5PfCOYxtViISxkh/YUpxNO46oS32BFkrvy5eq6e3TaJ9cuIq3Wxigy1tp6jIIIvBG83
CbBj/pvtAI3+FHR/uHqS1g3dwpOWv8t9NBeI+TCKCDKeAHRzEYsAk9DL0eNffc8pPgOEM9+ea8Qo
RjNorqMg8rX/cIom//NctOuWzf2cQoKehltX4d+M9ik+eUXonJjZTu5llIZNJMEdWIQu1KoaQBFK
wD5ZiicienB1OoeQfH7w//A9Gy3iWeO/jQZxiovSTQsHT5XDb9RfjDqzB9MarVIBO5q7xrdsrLeR
RJYziIR7lwPcCrGrNuFIsWoEA0Clq4rnhyPYQSQ/2RvO5kr9zFw8RgthRBJdxOMyoRqm0Zjcl76z
dhd3Ueuy6730mNDt2iKSmyl9+s9RGWL+6x55Dzjqy9sXs2QfyfXxiDiA4xiMJLJoaGFnmU+NAumO
x7glVTcv8UwZEG9AyZgRhDdzNnQ7nUfWxXehdOzNej7ZHGrKYN/beqUw8M+TcHnndoMyn7gsSiID
/1m71DNgaPnKPSxq/8nbV6cj7xhXAN1E7KzJWbJtTBsRukJ0gxo4MBYngkuuNzwBY/Wr7pps+gXG
c9OVbmmV9XNUZacoHTcc2jVx66cDOaADGm8yz5XHLpXTsw41nq9UwVHZaUO27MVMSr0uDH8956SR
5sE6kfb7/ubYPVRSQ4KHDcjKgXvI/H7QxbYEERuzpuQPTzPyuCDcUo+kKLXm3nkANc96dU4uraRG
UGavypC9EqTPHZ2NA5MNrOSSnOIFu8vkHRjh+rW/VVgIrHoGp0jqbtxyjI6AGW2WNCoFIQXsgVP/
3ti2TKoSOiZoABeb/jP6xsIfwRTmaQv0XpATXFFdTBI88+psVkPKY18DOQxljL+8GjF5LJnFBjtk
G08HCQrNwCyysRTN1ILefiH1WowPiTBXQoc5M5oQ6l49JuAONxhOlqGJrX+RkMcF9qtpCgiHJzxn
nmEvrr+1o8vYJCghbuDEjj0gsQ1PEDjZHztnoyio+dHcYr9BV9o0mM3NdBhf8kjj7RyJOhfn0iOw
5sGcT3tH1UJSUPhocCBB3UylwXLitAduUKafGc/2AiWJ9IAcX+8tyjyzqRUWDckHoDsG35Bw5NxN
BJmtHRL3lH2PMotIfsa+3Uz29eyUZNDemATEEf+U203RqeAjELwif3CSK4GytE+IHNr+jcW0nj7F
ktvhoNTfyBmZTcN2ZvX3LEbc8yD2kiO1RKsD3hsbvS8phIr6gxeaX+T61viY/Dj2mYn7k32+4wHT
dw0F1BHWoFE2PM7uQQqZYCTJwYXZh4SdW5rO/RvY5ganmHAJ/LgDN1I7Irqlzu/yNfpvbMcGD33N
30gpttrjP7/fEuAaH/Ng5vlM2PyprGoEMsZUay4zRub8tXCX8AabiAvh2syhOzgWnRJ6ZKgLnCgm
t12WImZavz03rmRkw4tu8KEDoBXfDdr3hiX1D70yZZVed1yE300VCEAeYNuMesTbqo4HJ6BwYb6a
Bn6Mxh/zuZ1uGdQOcU6Zw3+2fk2H4aDVkcDom6/ZdN1cqR1if4bh7NDfhhG4v4H6/KCCKqWj1ELz
LRdRBmHWernDD37+fYGWifEgwMp3hBaOMlqFJSwGzwloJLIT2X/47nqHlozel4zr5iTQV4cKUmsc
0SDzxzDnGUYpB0HI2HOYvU533cw+q6Cs6QcuR6xE+LKbHSLXxItzbAbdhRrjaBJ/Q6WqmtiP2KOx
xtfHoA7+XA6F/5POPVzvhyAmg18gR9BQq9VMWShJmeZq/nWMKwtxkRrF+Mtu7jH5yN3LPxJs4ScK
u7zXv8R9t3dQk4fFC1uosSSQitds4RNh1Au9Q8wJT0BoRPhLYpVguU9GnjeM6eD9ShErCIhIss5s
K8/NLhzFg16KO+fquQo2h0X9HsuZqD2KFgQI3EdTW8cl4t6VwA9VjDuKJ8PQcYDftP1BMiHvfJo7
8stoDnCjrjWIppJoO1wybYU7OGpQ/sg+w43xhN0hrnzTnXOamHNBmJDHkXYpQvaZazPIfBUt1CWq
A0G+NFd3EaOFNy5oCcmeeW4MO4QSDbuUK2DqWJBFgh09AvqwMdcU4aUJEfq4C2IFjdc0s8FxyEM9
8H5jsthm7qnYysCuXnPNGofioasPbtOZtQutDi19c65w8Uzzmc6TWwS8lBuLbFDXYIOBM7XWE9TI
GZ8ZG+htJsyp2L7MCvX6t1GlgJJBa8vxWI4/eYpJN067U1JiTYzeAX5097lQysgS/Gs8OJtpNevQ
Z/BxW4P1NOCST2huUiW52dFTlHejyikZu9P+I3UmcODQAJdtfD3Hv9mhO+13kg7WGWFjNuLBTRAl
SOIWdhUFQ0iQOn2NOZ+oDEVcrgqObeCDjFnyMoK+JTr7Os5rmMUt6o7i+uzECOstuf6WndUTX1eg
3tdDelNPCHFLoAw0g2Eg0KyZ/n0eJ+ahWg+PpnrMpnd50o1Y4gTCt5HVRYGCuo0CPKfQGIUlUgnV
XI1GQE+c1D68KIOAQFDTlTjkcvlL7YKGpRJd6pP0+uTluHBFr15rEX6TRT9x+fLGmj1DAQVZJLrz
MsM6cqs001Hd5FpIeDgd+87bmh4pcfC0zBkum5SJDHDFwWv3cCblqvB+IB5/pEmsnzJFEtKNe9HY
Zg+wLvnDjqNbI/i7ThNQ4yyB2iEyvmjW5VQgQm3AkkSyOaKAVA52+Dlpn35QnZEM873C/tGDGSKZ
GKz5LmvHwU8+Y0QsyG/a4Tj3W9uUip1mxuQv8EXf/3CbB5ZHDrM5xed5CopwZIztiVebvfg8faay
x00pu5tvbUxCIadWVMiK1JsU2wZUe2DzScnVoywMFGWkWrV7VW8takgsuENw9dGDTDlapiXW9lAR
8DSWq/hRXdArTNuMQ8uO40JuQAAW7DqS2juH3r7d/xMsWIopBvsstFKziZXhL9beQHMfIPb3CeMe
fINf076AVBycvu06Lm1o94V8iLOsgpaympdXDrni0RKH94eKOPzwkR7v9uyUEe3h5RjnJpNgShA5
v0cJqpVhfuDBBnF5yih46EaJsoxPEglFd5dnSkrEFqZJhE69jocvfyCrdIJUfJ47K7gzxrslNHtb
B9Lt4gnb5x2hVAaVyACeXU4FpZm6DUwnH3g6lLxmMjE5r8IixnI4m6hqQXpL+m6sfSDG7De+R1xV
IWBx4Qyx/kwHi4vGW9n5hBQTmp0JiehTrqsQBP4W/ISTR+MffQXN/HOPXMbP+7F4LfHa1jXJaBZ5
lQnlLcHdCL/cOmLi64Wq15g3WAkcmwsqqHG8boBjSbyl0ZIiUVpFrFSUk3envLcR0zsqFCeNtYkb
QsRilDIiKsUwB6+E13f7ctp1EaETOXB8N6f6M/ldJvY6SsZRt7tgW1qCp56SLCBv4qHnq4FJVZzg
4xFO9vB3QKi1oryMu6jTTF4APU0sCHwu+G3YVAB8BBcz+Jd0rG3lFYFM6vM3lK+g1UOdLT3lY2Wb
oaglEKN2G4z3P7CwJdzNhRiK0O9QvhrMAr1YT9r7cf2SjiqR7iJe2Iw6xv5OmW+pOtzPXS6hOMW4
ePmX8ieCbjLPwiFzPWTEnp+onUZt7ThE1XxDoz2M6iLPJ19H4jDBo9xMAD4UUd0mNR4rCsgxutjH
nn8laavjzVPw+oagDujYsjQ/L+78LruipMFnuZTEqG3/RnMexCryjFwqUKADM0HxZk8JoxXekFGY
nffplC6lxiLxmENPqQnfVtwx2KDzftJtd/k/Vtu42A+CZNzP89mgqgtg++2soH64XHY9asbWydiC
AlwW1QioW3GgdGdJZhYhUaxuLNqsO8qAOFf5F7Q3znTgQWrkpgmRA0M4GUOQf8u4xoommM7xZePy
WIfq4/b2a7h15CATydimUG3mX9gsvfoH0C2RFI3ZVWkLf6jeMe32qsiiSiIixNDS6PF23UwdKfvA
tj8PbbuRQnp2AZ3uciATiDK7lxGEBRqPQKJchwkbjFMOnDUP09jGECB2yccbPIcjfNhdHWLtHZb1
24c/YGrHpnJk/gON4aXjW+J4aTEESqjntrQJYWO/KU2naYyJO+eShjkKL3utBeafNr6vkaAFuxyQ
H+jze1EL0G5Qu5SOwp7wdq07xjjmys/jED+eDwp/sh2oiVLpSryFkecuTVTm4+2GmUmax2bho9Wn
W2k9gPcbwmFNLnBaQPoksKZWqfnGGztG9vkC4NJpawPMygfJsz9EYpsu8vnAERJ/KPoKSEJaDEup
BsfcT+n3sOl+9r5J1vWZSILHOxIw7o3K6ZtzCzppDwWKkDXYOpib7oMWr5YhwB/MvQMb+jH8wLVk
Xg2Ssg4ZW3rQN2MHCY/eINLbFqwoaZ/F7cgJHY/BZqvPb/svSR8SpYXRHtdo1E2kALOoTAU2s+6q
rpXRG02+rWzd97YEgvniNeBeySpkdFkoXihVKbbwWEW6twonfHwHuJIUXxoSQm1GEjqSI98Ppkvv
Agywj+CgjXC13X701afinYB4iVB1G3Cl7XiHFGfKSKg53Tb8v7SawJNdJiPAiWrYXw0lspMPNsVs
29xF4otivShiPLM4Fw3U0r0TkWnTOHIiDa4SXy6vgDAj30A4Xc6xNg63HneFpynbKwijhcV61/XQ
pDXWS0DL+r/1aTiaZoxZgmbsg4Wn0ZcpIiwBF4Js80AcaEkl/cCSrWToGxvQrOn+/nCYnQjiRHkI
dr9PBDG5EGY/+gnymy7hBbfMqqTPNriMm8UHDif5lVO1BE1yUJXHSgjlk0EuE5+0ak1PV7gD6lyH
csWiz5kzoBDYDl7DQyGTYBKa/rKmkDisf+zX2oJf3g/liDN7fRrPNfEvKLBJAwGT5rlvIPHRQBdX
HfVv8dIicJu6Yj/K8mZTMQXQ//nApSOtiP0wbPvbJIy6nUkDfSs1DK9OeNaPLAukVTYsOWYnwrGq
4P3kpMDf/wl1x01gg+CJ8mv3yRejPtTv3u0w/dSolCbnmQv72WjhQtsmtvykw+dpTx/iOXuSvSjT
QHDy7+dXWLLV0SG2WVVWYprLjNSwOTEkjBNn6coFSiqYNwF0naXtZhChBd0BiH7di6j9sz6+DuoR
JrLjyAIJUmXxIauqxvJmSloH1l0hhxqN0aAH9AUgFSBm9UsOrAqcFb6sJiIExK+EbCtK2Mtcs+Xe
brStHENimpTmwC2gBJqXhUzhN4Kgbk2DaUtT34wIgXhGDB9c47CHL3l0SKOr2Y+0dESyxRdzlYy7
sX6F/LTQr38sxlvLgLEpnWNRyvcfdUBnETKWKDfSp7gxIb6J6a9VKibUePHjgPssDOXYvO2biD+t
us/tDkE89nWJcfrtt1etMcEuojRZoslS7cSQGfv/trYKd0ElRLUsg7//6FxwOoYL82sdkplU1Xte
g1ZGVSHEBA8aUDWA+HrlQFApvlXHC2HDceTJ45LgVlMguyXpBbYLthqcLD6FL2o6eQHX/TW95X/+
QIjoSMpsQlKjhADgqvcXLe9t/qWcpa4lCToGOcqKh+u8HnseNOdWHQL1Ix43/IO0Nc/oEfd5F7Ud
2LE7NOQqvK0yF3OlAKfA1R9drMiHK60uTby+GIxX8nt4tupzKLlBgPWas6RzratK1HxGUOzEpQXM
0777cuR3t82NsC9P22LzxfD/8+QZamBuekAsIOejTLKtjFqQKvhaXUg0zuwtlg0XR1WMvIjSi+cM
njePvinGW1JWvHe52YbmoGNwUz/4EUo7aVnb65eZGbJFOqZ9f17Z4Ivd7sRgVoMMas9IilNUr2Vl
xPP37Rc9kK74KksLS0EjjvdDac/D+DtIq3yh44GGJdFREfDKiQ51QM5HEFVl/q0sESxQl8jp6IEe
SVuyaD09Bb0SyUotDfGqVMpDIfkaoSEFsdQD1Gm8/6xWx6udB87uYx83bWFoTKrvqbGXGh1SqiL/
5rhFYDTs0HLsTnQyMSZ+UycCqr4RNCZbdiBDr99kBoxNNdcHtKUZzajCNgWmLgTJ3/YKXOPjcbMV
aV2XN/py6vEkKDSG3wXXq+gs8MyyJvPZOZ5hzQjE8f53/GBx9yBZLgHWn1tTcXh6ujxX3s446EV9
/PUUK+Pp8+Ng8Kg46UknE810BS5KZW7ixJlC0/6KSckd5AmZ8M08EzCauHV+M2mbn1fxiGfK5P/7
GtACSqd/hwa2ZboXnj2DQfHCwkC99vGP+XRFFClGsZnSjag+HZ/hkj1OtuXW/C1EtzY0Gi3Njsdy
Nrw01Qeex3f6jvNkrM5aiG4iM0ftpKoYmI2PZHELrDA9TLalKIXEwA/bkrahbgBh42uyyxwQVS1L
81C5faN6S/J5FBW5zLDwBMzPDaLTMHxkCbmtI4qea07wtVhhFHpehE2EwrwZauARKqm5/S8QFyIe
k5X7c5JDtTqdE95bE9xHup1+z/0XmqU/PxS6WlCYNMApXp0iD6mjzxKYV5FStk6ST1U9UI30kjI5
KJmsr02THtruHP5iMo2pCXpdqXIJGKINPeVk2c7ZPErXgMe7Mi9K7bLghr3im/VBdm7l4SjkZop5
zRt7jJRTn4sUSPy+iYvhJ87MECAV6H/ALgC52Ov3XWjNiz3hVHRYQYC6SWbCAdJrQgacTHNZI9fg
yTCc1e7VqZJrpkepRdFJ/lwcXhEd6qkvJrt0tFmEklmbIvBFOaStnBIGpMOAtk8XJttIBcuv/Bxv
SmTawH5yGT9Ky4m84JJO/0VaRErijXY1YX0mAR6BjyloOr0eAs1iCBUgUB5DJAsPzPhGzqlBXQYq
aakIWWKRw08vyyTPD/xto086qUmpMLi2HbyAM3uHHyI17diM2yogWdY54CKWIHC6miYQyX4GVf7F
SGhL1oh2iXHPjVLL0MjTgZ2GjCOsWruyU2AvY70hOB3LddqVJaijiQXwxJPRdkAY+Vw/+DwS4JIM
3l75NFEwhdoI4yr1Oxxh2/7yT22t3074Gsxev/jjPHJ76Kaw6lxeHxsoaL8smpBVZO0kTCJgtGQh
oK4mPfN+/8dDZldxeLPr4Yef5vIHn+Svs22mzLh4hIBYJ0xJY6mGc0DXVaQLXtDcWEv2QJKrHMsv
sMTw3k/wTeTEctjf0NifaK06qJBr9Yax4Qk0NBx/IdYXb1KEdY3keBbi5lO/ImpNL81mLHP5LPYy
GbHMWEX+YOGeXIua0BRxml6NDKFXeC7iNMwtZPpt3SyD4xToDp2egjXUSWLU65zANxrK2MYyIbJ8
2eMP4cNaVN/Q6ERPEzjOZR+sUPUB65YhtN4Lxu0BcvT3SYHlPzvCch0cSEtzMSkKYN6zt/6vfnV1
/ksLJFwXsD/rih6VgGScgcfEBUJQB/iSPLoIfDJewPEGcyoaqDmpyNxhcUh7D3IqPVO6+iOyeF6d
uRAG9uYJ+V15cCPgrFILp/u2H6rIQsdcLwVjEMe/bM8VBqUUgqP4ljy4YHvDT6xWrSTtkFvBT89A
CjQY85HMcda75AFWpwmzJuzctS6l8R0e8pwioEvOk8Nr969pF9Oa0ddQ0tL6WUUJG0uNFu0V1FGO
fSd7aooM8JMpYOPsDbCoA321EQskCFcVgkMD5httzuvIPXwQPYofDb93fgO0rQe44IaVhMV+skut
5AwCMd9EjJlU+BHh8tqcGRP5KvhJG5zywSZnraZJMkPkb0fEg6MMGgLvQ/p3d8BenFl9BWTWbKkG
OCrrjYsJG7oZxPLxSqI0cc+cfXAzmICuDdgGpkNIaFGpJsTqO40jPxFv2cHviT28qrVgK8F1iV+L
q60hQxEyXVnwGWfXH3JfIUjFMggNvLGJqn9H7U3eWqpsr2lEq3hn/De7wKNvVRVE8IO4ahSyVpM3
ZHhbsnAnW6m/fSU4p3Xc2NmP7GpBU9FqxUET6pSFHWS2H+T9lN24s+IETdRagER2E2iK8eD9/Wta
qrZDLNOyOQEkyMxCJLwepxxK5zM2vAoi3WPfYtjFSex6S9MSGSw89CqktHSGnIquJDlwxck4kclB
L1hcMPeC3z99B+XAiXdpXk1OXRvgZuDEiK8WvJpS6tC7wiSd9JVnioyJIyKWBdr2pOajwUrD56SF
PFhyHcfHsmGUDMr7J528kxdBVLIgvW0ZWoUTjn0w6+EMMFm14KBDguUep1MHTZSMa3+ChaNYE4lz
SEar0d7KvA0nuYQSL1u7wyay6Zl1vqqiRDxBdfc/32dAD3Zp3Y1/0W+CKNTSUrBW0aI2VFjUrjua
xseJ+CxOv3a1PHo3jQjEjCVrrMrR/9/BWZ1ydr6sq1AvogkaLpROxgw8Ip7g+ullDxNmaYbxTCwa
JWAI/6NQUQp3EOABWVodfBZECMo2Owy3ikBJEHLBRwPNvcjM5bb9nuniI99Y+Rr/EXTNpcCSKXlu
Qtkhc56xn1naHdTmmcpLH7fNMx1XqKysFhGTNnBvakJjgcRpChxyGs1J6MF8e3KfgD+aP/f+ulME
zHqDIYBZLFQVqeJLp1ItvO0v+/HhYC3m3N1rTZ2WUQpjNwG2mpSZYCUNkEWQmCJ36ui9U+X1IxUa
yO9xBZdkP/Q/tjybSnm9kZk4W3PSkxszR9nJAkV7upUOBJCQ08WWsfoK2wD6mF+IwgBA9zu0if6i
+ckAFsRqr4Too3a10CwYhNYh8bJ0+MivpYkr9sC7ZM0PwwfsDUZmB3cCUghroCw+1kdLHZH6s6HS
G9775WCWifsv9pxO68SOVuFwHkJQ41b9ZesjcYDPyMVNIqZfkT3rxVoYvCZ+y8HJR/vGVz1F3Mdz
TsVUDjjrLAfoa+GbYGx4PkRgzseksx8OqmVVTPIWDacM/9L3mIHyag4B92xwdVYXPjMIXqw/RFUR
w0cyNB+bLjTNTuWcwZ43Axl2/w9zqKFHnbGj0UzjbJC8S2+HYk35aFE8KYe3HikpWMn7Ey+M6D02
+11hM0TFZJ6nvB5ufn1KttyjwI4hPItPs6Jq0F+rqnm79Sac5fkpBOjrU3v2yFlw5suRTHGoecJ2
dzKLbVkv6e/XGGNxnqSmhgyv2ye9A24evKFRnjyqDF02s88fi1Z+pVmznaFr5kkaiAnEDTwkXB8/
AgAHZOsMyz6Kp4FZ/KlyrW1B2wiRqpp/aRc4GJQroPwIB55+b0GzFaoCyEukqntwcSJ1sNCoklKG
7SQVg//iXs11M3hKkgMdWCHj0NrhytaJyM1Ol1aNGZY6eX/Afc8ma8fHoXaud1g0cq6apB94MxAL
GLH0QjxQ8MUQbbdpi2nti3NxSXuqv+SZ7TUWzsyJUcdmvPEE2995yQ5yvoDHkF+4N+6YuEllUUjF
xF0D851Cv37xjNn0Db6aNvwu9ljqUaaGQB1WXzYDmEKGV4cp9dDJ2OPCpDinBVUaoZtJ7mZfLUeF
RAEd6D1hgSord64LvsEFOMyIhnGqpXXVt069xwblfwRaE++Iol21fx/H9J9sFIgLI+FR2pZw1q1p
TAddJ16SJ0ugTyx5MJEWm5CHieVpcOEQDytBv5AfS6+/8CqqOi0/xs6Kv7IUA7D39p90vcMv+qfU
XqK5aF/vlXKRU41J/JJKkwyJmY9ZGoHv2KfO8I+eqIgu6hVSpQ0QArdQEqev4DuPk5bvNrrPEQBJ
zPWvJ4swuQzoyJuE0tg55nxsUyAu6jdihk0ksg5AqCUpLYxaxP4oBhi59PZwM0BFEy5ehd++4FCw
eNwNMeGstBrLR/gYe+i4Kk3tt3CpHhzZd5fdd5xfdsOHHMJQTM8kzWvHcMSLmlUxwgTfVqmtgFsa
/Crit61vMvx80MDuahFiy0apOV13dMpGSr2wS8zSdFxCyTKSf2YcU93mAxY7QBvhxvq8fEROEfQC
y634JOr68KeltH1NkWifs4b8cCf8Zq5bRLBHpAtuVVOd+VmDVZfZONgcuGaCZ4krFbk8hJaRWX9I
0V/kLTDjsclgXyFLpqXlVsmbYY6TCaB03sd0DZtQgs6N9n0FxMrzndthVu5nN8RpCMr5D+bo0PMU
4xT1uq910AAFdDucVegYdLlQNj5eKf9OamxtMlmIoLYjTGNqrTsf6BqA+Js6qFMWnXuyE97MBhYn
KP/RnxsXuC08GCJT/qCXjN7UTGIHZag+sOSD/GEfvrhLegzhn6D0uCdd0S6RsEHZi7IflEz8qSkM
ux+9rakE4i+gH3yZ2ccUjJf2Y/UTLGnB4P4+V/PHjzDzwsedAMRmLSWwNGfmSTUsecIfZY+dKrWN
q59iKBqd4BcLhRF1dqJ/93rxGtQ7/Eg60o8/FtvF4WoTbQ/DD5fxNcilwQH/0yVo2dNJ/IMyTuP6
i4sMNgb4v8a57vOn1luSn84lDNskv8JAM+gJbwfLG9j53kCIUayOZxM6u8RD3Wx0Za3PIpqlJQ2c
g7O4h7yMmsHuJF88FTQQ0EKiet2/jkgKvrheJyWVV6C4Z9Z/0itBlglY7O2q07dA/C/xTY0N+akl
IYK1aPn+4kwlKHEBor4pMyHVUFB83ljZdZ4CBDVxSjyt8D6Z7EDe+7jjr4acdSyiCWk0rFlTIzcP
PUtPwz5LyNiWH1+cN8671pSZuhnp28hYhnxz98OmM18T46ft7OgypcovUD0RmeNuSzTkbxehyFlb
fB1x1Ozz571xD0SgCpZ6QIUzQ2uIXTb14a0QG7DV2SXkFeMHoIwcdTpcJzk2vRKhjnkviI6GUKI4
ZVKs/nSl867bR8e2RTCQm1pvGECF+IkIWiexbOMnjhR1GiHe+WKgtXuHwC02t8CXkFoCrmWKGNdp
2nJ59HD2qr+5508qwVJiVEroJuNamPocHrRj3mVQFTJxuFi7qkj3Px54vz9CIeAUjz8HDIseWyMh
Wf+UL2kvQq5DOx4/dkIMQm+0GhvfB/da9l0/9tzWISnEdzKFZTy83nUW30lCEAbX1YEqOUHBCh4Q
NuQtgd/fWgeXQjkFxZYqlOFPRUT1hJpB3Rndnc2CFeIU2cNIP3sZK98P7igPg/joviRuyKdPu0aA
ZDJ7L7kDtzD2b4OFlAp0qv9XjmjJthedihcYDItzp1wUw7TtX9JEedGZ6ebDv6dHG+0bYs+7Re6v
FuUyg7ptfn7KquqqIa0QTrz50DWWk4uibd1LnQxgBodLMxkI++rYJ4NwWiJwXANAyGhUpycMqffJ
dUR8MdJA9R2TgqH3YT/I1+RGbwaFTfGrmfhnelypCti56CM7BT5IR3SaK2k8i5KZNFy5rFlHplia
S5aOHDFMxkPZlzlDYM3oRF8GU2HeM5OtZNSjyRClI9Hc8sXGfd0fr71tST9+8xZyVq50N5OtSP4X
/D6kDWTpnx+a3ff/5Jhmalmu4axF+ras5NQeGL8I7D4HWQLQqcF9AXd0xJ6HBHeTguihxd2d7St3
iuywGecgmf2uRPKykDDnwPOBn9mgYqVz8Yufa7ZKJBEbQ+c2Ycxl034shHwtFD09959migXJ3Jzt
XGRf2/XoR92tbvucBRJ7S9GFfInIr4yP5IfFm6oLTsBxHtU1aOCTOTcFkbOnJivGW4DtqEVGTCkN
GHSPy2GDQJfmLp4WvRmA2kUhhNPkz/MrUKZcU9NA0fq16Vna+5sfRwbhFqnj61RHhcfsOEYFQM17
JIeAZw3MNUGo4hkGXjAeqhYVSPBP27GueL64bpAPaMz5PLCU2iinBVnx34MCN8veLmDiveyuTmwm
nbHMQPn8sm6KldQfbX+nf67HzU+GSIK/o2bX79Wevwag1KzpkepNfpC4d8ghYhnETN1U4wOOCZTM
hko5K+txpsoVFxVWz2JOa9lQ+yaKSVvFSJQeP4dDeW46EEuCNUcA4SCbE3471/UPFub1VhrsptHb
Fy/lExxGtMXVii4igJOZR6v8FqgJ4F3bBNvicRGwPZ12NRA1FWlqXxgKr/IMspiuBNd7Unz4pd8a
bm9FWOvs/jP7lVvRrJs3ynvK9gs8/qTLzuBw/BktLK+Qt7XkeGL83LXFWCr7u+mrzQxjyvos+e4c
qwVqw/tiP4OsNq86h7vW+dXtNfbnPbBf5uo+k53JU36x50FzBbggFnNYcR+3eRicjDyM3iTQtMSG
3TZtA2IRcoI4I/UFpAraZDHN7wcqaL40ustgq2QkGkJJl4caNMCR9m8gm8gEVpiFW36nROI64IYl
xcfzmqdu6vx7exUXZ+bnxLx5i5Hj/5/FmfFBex1bm+OD5ybZ5C2I4Q2xtHyrNs+wWwCDAQk5wXnU
iNBp8D4BLymW1fFIQowJ58pGCHzNhPFP3aAnL6/7TQpIEaD0cIKrSaeg4LI9Nkr50VeqPIpqBSrS
HoJ29ZMbxY7KiOuthUDIewrqati4wTH79aUgkaSU8Ho3Uy9RNW+RQDiErVKcrK340KwxBe2hZiGv
XP2PlqAoXGnvO0PbqxUQGkj7rmT08wiUuWW5LxNx3Xng3n8Pp4EoAqiLm/Wj6JUbixMm5JLlecYU
C6jiuH/1hnDOCGvs8TOa8PILiOEP6jJzvzYsAyqhb7UwLfjDvDVp/P6tu4l4LPA0BjNsokiK+ZYQ
TuAKUdZLWDY0JvrkPsXsy2Oo/X44/HOJMfSsScc0xMbQYSbUJZkdnVjDaK9KQx+n7pqADkD1tq1W
0Vi1sEFZp6GQGT7oP0EbDQmgpNy3iWvIXjwvJsFJrCuslPelg1Sp8dXFTPcX1UYhD3K+ZAUwUX4+
uRsyryLyCmLSojCh0OSp1mWK43TvNVGO4j2cKDhUJ15pK5jqfAeDMwX6sMC5L0BLfO1Qs2+OxPiW
QmsUefHnoAEFG3WoQL6/H5boXUVnmFx1pEWZoFzhZ0B4PI9t+Iim+TsOmKV8+bb5O68izkFwXDbj
wxM6gPE2nCP7uuHDRDP47Tal9ki0FsD1iUlxE5EAaurfffbT4V5wt0P5YTfWidxf+Fyp6Qb+2lj0
dQm2zcTZu+bSx8Lx7hPcqkRJ1lhjQvTsH1H0XZnRQQ9tvay7uhfY5muHBYVRUcmsyhAokooffv+x
xPIdtDH3/82paydrFWHRofR8tpuiTwtmHMfzNLnvemiQi0j5gH2XJGjCUlYqKm5pv9ithO3CGr+m
H19lPu7eAEiCrDCa6yaRbwqihJMBYlhDOu+pIkev/il9YTmOof9hbb0OAUdGg8zr3UE0bMZijti+
2hX8L/bUgE6F7M6jt474cXfeWBB1A8/7OP/8hGGlVccP3AeVIHVe3VV6qMkHENoDTnCc4yv/ZWdw
Jpf+aIIDyQC7MlHHzUNil0OVojpmjBEmnTyTxrS+/gU9N7nJenVq/HqxVqPM9oXTUSEzbfi+T/ao
IfD0jlB6etHeniZSuwMbJ+WOu9dEQXU8POrra+XrvaozTp53q7C+DOY3kA8k9+FPJcXL7NIPoUeL
e2NqBb2IA9pesfV03No7drFsOpmObnlHWg/KfawgWhC+lt2wth9utj+VuYILtbafBnECkB4ykgOj
nUxd691kUNOdoxAV6kKn4i0Z74X1k4jqiDJpSYwXZUuWEVVAmrqa8MZk5MTA+woldB9edeeRtpsS
HLvn7vcPNIyLKEVSJYCuElbD2aWacQZ+Hm5uqMUVpDl4rfeg09BgLBtk9/7ErA6PF0RUq2DpUUrN
stZQ6+HLnN+18QQwmdA0JVVlw4+/YErn30thste0nUCONJYhD1MLUuf9cq1fzLHdBTJblIOv92aj
Id9U/6vcVkqicu095vpaB5rQDtYEa9OJzZATwfGzyi6tbkJ6FM5ej7LTS7nklj4oj/pPCs2zqlnP
viXMhfCIUOEpTQlPrIsVxoX+2FQZ6az3FfY9RMID6NiT1gZYOkniILudmRIo4UZYvesH/g3UPFlM
ktiscctA8tctS7A4cngiQ7+154GgZI3KdJgw4jhasJTG8YdTrJOuGGAsHTcGbfhf3gzwm+mcMAbd
cKtERvkvMDC9txqeI6fAVV2ATriUJ/RPF+99wttLFPyDhWahVmUc3uwtJAiRz+C0XyqnTNSq1AkS
I4zCjuaZDSfk2Wgcs5Ghx7Ju9TO9wk8e42UEenPm634mCM7JPr0GTvTyGO0+Vtq2f2/6nv0vmK02
hX0AQwWI8cNSCEBaS4eBw+kGu4cbRMP3Kgd5MjH8RjfjeWCd7T3dVenHtRxrGSzY7wc7FRBxzbSm
lGx3qQdvHtkQTVoLwKVp/FvOtPQdVgPDyWgPRvwACF/wKb9nUiNPGOprNRkgXrUIjplDD880nJiQ
MyKwvfrVH0NZfb7QCgBqT/XG5ULozWzWir8gFRivpBGK6rOLlVWXCs+o94uMA5lCN8GzQLNUinyr
lYalCT5wpd9fsE6CqyD+tiOKwNBg4VcuLVAbb3AIwhmb8wzjRGujohm9L/D3FSA5pisQD82R5y65
95ZWJxiYh8xxN0ZSrYhE9aPSC2gJsg4qxo28B5hf0TTeqHp/JOd8y7I9pJPorcBEcBheqTnFNS8d
wVxEifYm8u67IyDu0y3KUU3ZUaDG78FPPpSr+taIjSLmX+mpuExqLC2dYrUem0nAMRfWppxqquwA
6lqocCUL3YOjZmiEugoaZ/dnI/bKBBZiPHNV0GSN0jtqpHKFuK7elnbsDH3DJMQwS8CCDOrti04s
pJY86fDJW4k2O4UTfAT3oceHe698FDkzBB415zq2IYBm0Q8oSa7dvOMEhG9/qFiCb4emFMJCEhX4
ZP5qGJwDvON2a4WpvK5MkYdFQCFlPfg91dNYdADROm572EXf6pcsD7fPlRpw/duGJEj9j0StmKOH
NDin6qmN2zPAwkHOrRystqYDda3FxVnbLWypvSMDDZDzD7jn4XXHvaNxJVOnRr4sigVUpnY1k2zE
BeMM/zwl0mAIweDhpaYwap0wr4shRDMS/cNWii1U0nEKIpZzGeD5l5zqqDZJ91O+IliIax7U/qWX
aVSCOHVKa1aUnOl1GOHPNa6fRsTbQWwH8jxfKfc520Qf2zxaMpZwm/GHE6B/v3hWVmMld1Il/Lrq
PhIBPfkBWy9V0z85yv11BA5SEUu8sIqZM1dLSqoNyLgfXV3eiKmxBjwVPILQyQhSWo08hqR80dZX
5Ec/c8ayVifALqL3nA4meEE6qyF1tbxoRreeDcgILd3qwKXurAH8RSOpA+29dQTP+5jgbBNCqnq7
VO5HSzTOe5Rq/CbcDYjn1K74mSEyJPP6Sk/Cs6iVT6RL6NJdZ9mB7gFLn/HTVHG3MAJ7ydNkWSvg
/BMxa03LWeNsSypS01eQI7CFRZaPIcGoCuD8v+8gp7orkMo+6yQMHiLTAk+brThSrF2YbGR4Eq7U
6h5PaAASpa48MJ6MA6U4S61IyJdFb4W5CwsXBGZ4ZKzrggFTKxbLM/aQF8iLI3yew5sZ3smNLLLD
FIWTfcOEJiyfkBfVwzSeJ0oOk5xrcbjuslXIXmiIarzgqDSLNiqN8iWa7tgYNaLSbEHKKD5jxALU
H7hrsyW/PUAktihamOb+oZsg6EaoV1S/w7MXUjxpKfJOpo7/xto2gYL/qD0TwfIGHX06o1Kkp3I8
2yrasmqyItG9m91IROIeXHJTFzOlAGukPmm9XYA0vBFrKD05tjLYMikj9Is7yN31PPw48np9JudP
L0mugo/73FAm+eU3B69LkAnAi/L2Im0cEt4U71hL3iYdd1+J34dKTESn26ZkXMxkXdI0iSNlpZCA
DNoQOqr4BbAW6pofWLe71gHJ9fXulybvmb5SLcfonZDpOomJ+K/pY5/jaJ1r3Sqi3ZqxHHSL6t5v
FNmG/Dm/Ly6cDG47Xww8CbB470szv4y9GNy/m+QzWy/8cfTmsv8elso7pDQFgVSyzeNZczL9I5SH
xEJxTf63Lb4rQvzRiZQovnWiPuaGOJQzN3kQX5dAniildR5y+dc9l8ZjvHecI23t7GOOShbSiABZ
NCn7beuRMof9f0fr5MDeGIQJnUiv8hyLp56gN5Tjz2R4+2nF+5rdyQWOoT0/LvYXyTdUt3nzKVk7
knN55UtGotns56sF5syFX3ewpajDoc/NfuV3LWqSbuEOb6/Y0Q1AyAA4iQmdTVlTaPXVPtbUBitD
JGuld+xewjjA/O07Uvi9VDt05dgvMB+uncVSC3WLrULhsylmp0yDgWlvAVscvRpPyWiWg34IKEog
6CfZpAxjWi7Uw84FA8l6aYKul5OD6ON5Cnt8oUJfiH2eZ9AiRgJpbhVAdqAABptgoHxBd9pkLLdX
SfB44PwZ9Ywi1dVwb/6xLqn2MVXdZK1JskFAp9aIdHl6Ctjc3KWEnYK7sM37jQO23MvQnVXC6+cu
5/uBgRCo1nuhlk5MBkxPiYsVnw6fF30DRHu7KQgCxGqMEfRfABgIIwUWpRA1V6gDZkc7ZlTFQmQb
v2hoGYf/f7OMcQhmtVjbY6i1OJGe3isik/+cEi9jjtYdnY9lIjCza+jSudqwpog7sOjtVlraGkQo
VQ3NYwt57g2EvKgi8OMyEb9q0UIkoahuHqDPkmsssndWET25Dai6F09cZBcDNlIQSkMERLfJwRWs
YUhHHLEDUj8sFQhIEA7kpGic8Xt2Xp/iDun0V/Sxf7FTiVhqz1vyeIhzbBNHCvcquoXFOcY/GvgL
aMF9UCzUA4F7aMNP3oisGN29mAVW+vpLgAWLDugTWWFPeb7bZbyD2Gok8DWGd3ylpk0fKSLLG//7
cdpb3sYvM7bb1jVOmvp6/57vK6X4ihnxlo29WamqqbCG+5KH3GtvR6WLT/dPb4B724a+FGQ8IaFh
jS+86758DKwo7bvvZS7RrajwHOG+XXgQJ9EIS6g25ynC7uuk6Yb3DTKn4t3v2+QiyM/iHrubQ7NX
Gptg8ffbhdEz4Z8zlxl/V1BLCBz2xKs1GoqgVv5oKhKfjZKWUFH0oku+w3mjd9tozUKXInVb2Ua9
EtJRHVVTGuju0URWjT/GB/jxlCXEQwkbLC1pEvHpq5jxVEWE8nevKeXVP07P9+Oy7gQDeS6bBkzW
rk548GHjFSShpgHK19QtRVIq4swGP/lo3Ir0nffpNQESIXrn6cxY11nRT7/3F0LRYPknFGBTrm6R
B5jAFSTGcGUkoS8eADfMWT16HI6OiZfWl3RYc+OF4L3/cC+b1Av8umMSIkU1muPhFfzADo9Jo3tZ
AspL1mXqnxXd1scAvX6V+CKqwJSI5CJtzICx+k5To+RBXH3KHwfrRP2fgDzZz4ZsgSKvoVdp3fva
fHCbsSQSSTWJDMOmxZe99HhLzzTL1ptWFmw57EcMtcR4l8rFb2D+4eEUlCcDYvhsvvG6wW9mYW1q
V0wceRew23X7PWMgqysjsF0HztXkzyeBZmdD4l2l0EtSRpfz8Zx71QvnNiYSW66Y5DhMEs4l//4A
f6lvjz4a/r/rIj3om0wsaoipTVuevyWlj6nEiQCFMV4E2CmYfM0ZqkMjrBFNavGtphCaZsvPfsMt
D0khh5zOcjFjxhXzFaqpbm6I8A/vGjX6w2C1wERXEw4tG5YMxS0MqZKasKpmkqTkuAkXlWWte6ne
zixgcweLXMckVj2RNPrUtB7bYtYOrE5dB18VQUkmkmxNVFQ9dZ8L3wa5F5puzQ2Odc1DRDXpGUgE
sMK1SvFD0+Igz4w8BNLY7Ua2XuRfR5jCudHeRgLhp/GDw/ChjggJ8u7CqMf6mTRzwCjUBQDjaygV
OAO5uj7RHoymAGNBwGjDzl1jtvBaX+v/5k79T6cdnVJTNb0J+XuvsoT4ssEPUERCqKhorrkRJv/Z
vQOcDO8L9xLDG/R6b/XsfGGHh9iBaDO4Tub91PLGweBis6nvndyq2/i6tXGTXWo7spojWDEwrkoo
wltfzZCyEf3j2BLJVjhfuPLGrBAoI94IhmzS+4H4nmXbJnYGzBlThfleuJjQef52Yy3X75owQHvO
+VWxQ2ccyIXGth9pukxDClkuqkkg5jy8+ULK/taHWfp453gKZjeccWENcZp0I+feSY07NS/3RXlL
894dTINu0zunUAQQY5tJf8srB9tg8wt5OL2C2TZRuZczJDLygr8QkDMcQrVl6UV+VEgAoLRRKIaH
xWcE6+kVmppFMR7y74gppOYJ4tWXmWDHJQXbzRf5arUjAKMneGeqdsRttQM5iL8fy5jU6JsiDLHB
Nx1xLqVfWt/t4pQzq+ywzL60C8pEvjawCypkqaJbqnSaxEqazhrZqI7UvT0PDhLcBKZOAU/JCS8B
OpotQPGH89P6+z5Ed85cnNtdcznWerGfv98jgfwaiuuwdMhEP89C4jB34SsVqKfmd/l/s96LUOoD
Rvc3POTYp42apc4+pA0PRPzMJXUA59MFzh9Yt6aJyXIOKPnFaz9Ca5jfBpldHFLzeI30JyYBrDr1
23dE8lcmP8HV+x2fV6JR+NVfwXCoyh8kWO0KNO5xE+dIv1XHLU/lLZJfsBRZRUF7c3KYJ45o/33j
uu3B26RPpTJ52lA01I2BrPeHSk0jG4zGonkBtIEAGmsrU48v1gOKIflZwn5z/LL4Byoaqab5/SvD
bJULFGNY7XYc5OCp87BHMYEqwcCqTRhK7ZdtFbhytfM0zmAzbxBMf+qiPRphDwKrlpi/SLaTjwCy
BcjBQ5XzNDVCkIG3eafeWQ4HhVKb8XN1kLP40R2V9OTYX/xTr5+V8gdvLLGK+Vwtwzs2JDkmfrUR
OjDDqRmqeHI9e6oi7fulgNKQDjgIlukRIbUwi8icBDScb5ZSFdtLfXmWRiFwRfAO6XzO1FY9uJAj
3CmFGgxZKtHpLMuCPS37US2TGmtuR6XRrfujwKrX6yxjc39yn6uzjMDj6sKGIWE5EkaGdD8o0niD
3z0w2M55VzUpSOlJoTxvsQj14+RF6Gz4TlvXkxC0NeN/8mCZb6f8X0cRK7F3m6p7/zB/G6T8pREu
2RlTVRLOx3/dW0S4JD0vc3CMdOvY/1+kqrkjWjh1Rcx+80WDmZD4VlEbZk/bPjZFmAX+U2glYykY
lwY2wKDFOSY7ovRyuwJpvrCMShHJIIBbYzmF7YJVi424FiwZRwuk1LnnFJOAnXXAMSFDdpxgI835
K/1kZ8pdqPZ2lPtygOfLd88LnhjAIuiU/piE/N3JlOOqv+Xxsnz0U1E5J4uRDXuBfrt5s1y2j1st
H+TwcfZoatSje4NHnFwk9uGBts/kPJzmLD6DZbHIIACxgwnD+IaMBPTA6F9ut1sNC4sKD7PgIvxk
idGiM24rzvJOYe1d8BYhwzMidcCVNIgdcab/8XbnP8k7EyqsJbkg3FoFAOMRdX8VNTQ4dvExlEl1
tZ76IIi64OturIrQOHQNB+uZliixYKH1AxYAhixvhRFdjcZUUi02zCsoGVwWvVpn2H1RasQskuBq
S7uph8U7spbgK2zJLX9v4RF9CbBtGLTK75uSPZu2F//FDFWLwuKilFfQT7G19CtUK/u77S6nCKmC
NGzEwfXxlQm6F0BeBXDkSBnOHl40mUCzTTabeBG7ll6KbM4U289SadULdOiEKbodZbAK7EknhUrx
HwNsQy42RnJAFQMCjXQASf0RyK6cm2mEhzt9iLHB7B+Rb++nH9oATgaXbX1F+PoJ0dG0Lz6q+gQI
Xq08EPIFKpPWByCR5VZC1ntmS8YI4R8WjokhJwCNAeiIv5NNECQ0MOo6/jCFVWKOnSYygl4cWuRV
LR0hQ6/LRrzTY0H0dyzQOuDYVa7agFPulXwyiHcoM4f9uQPKR7zDekN0SutsPoSTDD47lWjWbXME
SxQgtHtKyXdz/VQJwyddrz+9XMXCdsPriJfz2AJi58gSNG+xFixD3lHr33hnhGcll1G3ll5yxG0z
eY0LMFhVqcyJRWndCL4lJIH2L0X8YZYsFRmNHuZ5r+/SQZEUbtDzNb4bTfSFAZFnKRax59/XKkRM
8wzV7YJGsDIqsck+60BtLiu8Wa9NgvBHDySaIppZCayfKMZOdd3iaMugE/n7RTtzgYlg+LU6CxBc
PMxn6gl9GcSEecxIZNcKsssUd4GYpzLaCHB0rT3EEvDf4MjkCWE108exUONIJm4096KTP0lsZBGk
jN1bRlIVgagNOywnT0Beza21abfNJDmiX0uFApnPyGyTrRw7dBwkq0naADS6c7z3Tp5YT/nnEBhF
dnKrYCHhLlulk5+QwLp5aVMwoGTpn8KTC2JHs4YS0+oq0oJt+d8eO/ESaKS5VvaJqkdmF7qYk3qs
4Rpo3TKb+QxSekZ/LGe0tm9P/k1Ovhfqm/jtztXrh4pu+Kp4utLenlIHTKed9xBr79tu0+HbV1Ws
Oc7BDZNgN4mDn/xrlLiPM/ysea7hHO+zKOjP7HpgEKOPz5aVX7yWONe1qJ5qc6BzNngUIHLFvWQL
f1ZlSasht/WEC+ru/k5pUn1Wm/fdc3F/C3i6Zq9o95D42AMN3bv1i6wIOjlRK1MOzC5zxf13MzkN
vnt/a4yNTzkMoUrescblakKKF4WuAfni3U/Z4B/BnYW3E8ym65hgRn9jnQ0VyxJXgki42rBL3jf+
Gr2eyMghrSr8L+zCcOUE1mfN3Zy4hSq14rBtifyvRjqbU8YeuGkScvTaXED4Yv2hMfJ/ziwiqt4p
MHB/FyaL9syKg2oL70gGKTV/YrtjHU4SCHL0EBGZd6X2ze00OL08/OMXFj5gxzLDnHJNopNf+vi1
jjj5RXLZASCRQqJa7cOLJ8Kr76DroCDW7BNd+CLURWnOu2P2UUSTAM2Soa3hFf2+SuTPr6FJBEDI
ZmPw/aiFhI4YNfrmW87+L8SLECXyeLdN5Mq4xdX5h+dYFvkrvzcUEYk1+Ztvz1/JhQcURxm/bcBS
+jZabLiH4VTjc25KSd7/3DtMjKgykc7feESD2SkRgwO7jiqLlx16wU2SIHHSkJwaPU97YCluXntx
rh6zHr8akuvjPByNLncL0UL5JBZiQvZzQ/dw2Cq7KDBTHdHIpDKGSSozHp0Nqi7GeOVJA8gJOn0r
AI5jkXrrLfo0ET+rkyqdFArQxmswzAAc3je945j8TsyTLDOhKkxbAu21uA4ZCrIFdEZtoj60nN1m
z/jvz2p9+62FamgqIKH/8bJD1FhgIDsp1IDqv/Y5LM762xgFTlP6YAd/DRcNUNW/9+YCNn8TZ6IG
GdGAgnUnnGmDC5TrzqpqPxC/eO6k9Rq9saSRlqYX63+8HuUQ7qh0daCiPxASKxjALcePFdlQntT3
zIpUiv24UVAfYt6W7HKO0LnT2OSzCpifTp/0i5e0bVYBEEPmcOVjuQXU51BsHHNsxHiCZmwtETrK
tP5l2MoiERmOnL+UrAp3kqATsM2h0oApYxzprfx3zFNllRBpKWH4NrizAFejgClsOnhCW8bGhzoI
fgInjmgI8rMmCrsWhdYJHzr/yJMDohOKvYMq1587YBh6Xm6B0IP4HZEudLdGOhjmYxlFr6xirn/h
rqqyaVirBEJt33bAdqgGbAaCAs/b7ovZTozOnep+flhINjCLDdUak/Kz9wkL8YXA0yf89Cpp6a82
kXkxCN9YDhv2mxpyMiWPRiuGkvVLNAtpFTYu12wN/YDmGH90zth83T7w5qK/+d+C2uUN+coixJL4
R8iqegRBGR9hj371HAXFuDi57fhNjPBXuIg6EiKFiEJrHYKSD7NeTLvQuVci2OBsGM9qqs+mQnln
W/sZnJg3DMxhKbjOCMSFGBXXepXegRLkFidIKxXFojxqCc2qiX6gvqrwK4Llg5z43ekQOnd3zYNU
1MG7U6KnH8Rrt+DBhFiOX9ssiMbuSDTcvprWYcRHL2Kb8otfWplLGVnCrog4H4YlkZfOgu6r+jA8
Bywoy1vvB4H4eBkbIbOiU4GliIZW49IPPzpszDpWHaF6OwErOOsgsxWXEuvxoPh1ESNR+xJ2kkNR
V/w2/C002W8yDwlRLr7Fq1+A4Yf4RwtgvQkyfC4gt9ljfhBXE0o5Ilmyh0HYtsdur2PdInkHGec5
dheuF8267EiFEkzhIcF5hlw01D+Lg08tUMx93Fx5cpgFcWX0azVZfRnt4O93MnL+q0+Y0mx3iRuC
w63b9Lufie+6qdlNwomqnTwhBDNJXeNBKcFyoX7zkX80PWXl6cHT5UAUEH/hve/BKAiz2T0S/f/y
7gHBTuQ4atLY5Z+7SluH2fDGBmvObc7tjWii7cvvlI5ShnFprK/QdbFASfDjhn2cNnnnqrRlvQNX
8ganMWyS+IGG2l1S3cI2FmBKZU3lt4Fsh7KrTTLqhNPKlhV3dQppA34AHBCoEkiUzo3NScQWPZtM
HcS8BhchC80Rux5uTwU2OBY4vzNW0fUWqoUb1nKxh55nEtx9/KATUOTU3UIXdVmRu2HgBMFZNd3Y
yE8Cp6AIHozCrvG6p1woD1pgoM6MoL6W0BMQBkIZva2KgpwJZt8k8R55e5uFkZBxibNTGpiGepDS
xHzoX4J53m7HOnMWmkvLYEZ9ysiNqA2RkeVymDWrgtQGAZ42yDfGeHi8DFeF57YgIwpYeFs97NuO
+PoW6cVumqhU1kPBPZ4yeGMyf6uIEQISXXBw0iYpy/32fovgyHDejo6+o6wdAip1U29KMbbm5SrH
k8x6EToz9BrBpqanch8bEVE2HT1Fu1km0O3RiYyrmbXpVAJ5LH8gPd9RfJTRgUN+YjjysqzFZNOV
ggB08Sf0qPAAoZApKXxf8qskiVXAdAX5mMGx1So8Qmvywr/wjVmNegLcVL59RHKFjW1/BkHO62P2
/sHGoTPjgwyBSy7CICoh3UTnIEc9qmFfq96KBXeuK2qE4Pefcx/oJklGHmY3xAm+DidZGKr2sY/K
QDBZ2pNvcCzk8nAbxkNJw2ebAwDMNtCzw89FG+yK1m6LGsyCeH0lnMTTZnyTo5ppoh95tUIw9eui
EtvDyOKTJxi8kxy9oJR1CuOdfaOyxAldufcCXFvLxI20jKnd3E7WEOgmVKV1zfNIntZF8bK73Uko
hkSzyxJ+djL2ITtJkpMollT7BKdO6CDS4nOkGIDB9oRqKLonNT6W4nGIY+xquZuq1ad2sXkhotDw
BYxEjzCpznxYNv+VLBmkaLORHn4lAtJoALIXEEdVWxEGuoZz8qtGZDwD/nOwbefeP/NezB/C6jvi
0HDeT0PlkjKmQzQmxlCEOLV/KhCuHVGhOL5tdv7KJQwv1nFdFhe85HMDp+CNCidAPVFkJ/Y9cByY
lBOC92VXwv1Xc5FDSUzm597T8YOtcSo+lqhS5cppC/dmyAwDZRT7ALGIDsN0Jky506wyJi8ewUXY
FwNcIDlMYnfs1rh2YxApwVSgXrtAgBMsQYoO4NcLMx6iVX4TRLL72IFCq/Qo7PSurxJ/owlspYrB
ECssrQZd8PhafbyB/79IOQ2sFRT1Je+4BszlN+CUXM+HFymqU9oK4FDjTscQf0oTL3bbLBpldUvl
+gqOupqjWHLJbPkL4zVGWdwP0xX8+qGRC97HGj8GMopWKmRE/NsndDZAI0xoXxPz6U67mrFteU/n
qEtLiu+HqsLaNFgJNmWWaPtTqLD0vnHhp2U59VTR9d8VKm2WbLROiskZGc9BNG2/OvFeM6PYdKSS
JHkHVWAHX39LS1/YNSQCbsZ2sYjRgC8Dtk+8XvHfkaFDOKz8T6hxUDDhVuvVroVxpeATUagVrLE+
EnKvx7fyB7v9pKR07zMu1YM47N0XQWngoAdm2mSksahNIkjv5vfuSsBPaZLAKy8ar4GTgBHws4q+
QJpr66FKlBxc3mfY7Mh20hYncsJ62gvVrr0vYhpSEhpf9Eyk2i2C0MymWRrRElV+/HfiAMmhGCPL
AGqH8aq+Ak8zOWu2n4BfkWOJZnOXTlnsAtZdhllN4Db9pV0AAVtYALHtJjxziuwXmcMaoyfzieZ/
2JI8MPFdNBpgwEuP4xEdzKIO4OXFrwcjvfMEFVnNa02xx5sQjRsO+N70YhoQ9ezihBzbGMMJb++b
g5iIlCbkM0EbptnwlsUCvS+jPVdCEYwGGvIh4OSWBZxLvckuCBWEEGpFIbm32tge9s9dS8qYMDRA
XM2rQJIX8TwNuZtuQsHzB8EUo8XIwvunqcjdnPKGO16CYBuyXQ7glDRP8VFQNa1v57OBoc2YNF4f
xzWHHhDcpL1Chf9HQrQN8w3cldfyNE40LjEsAI6rBNJc+a2JTj1FB3VH/yqOxIquGkqwg2QEwtce
xq123GvuAMLTUe3NjqnxG7hKUgrbGwrMy4+OOU6V+Qhn9AfgbCADf3PoPZ+629SyoTvxoApGgyKm
4kiowIxrEZTwxIGcDUuV2KqOc+dQ0xm36T1SvC376sIaWf07QlnZV1TE9Bz/BNkl13W1duseP/oe
o/4c/cmZHYPJuB8Zt33GMRp00JOtmlXa9o4/CgvbMQ7Vc2taTo1gLYyoNlZXbfcvUaMXG9q90s8s
y0rNN9G+QXl2vl3opvk+Qy1Z0yS8dxDLqEvGCqiH7MocXqczoDiun4raClmAiZgHnvlozCIh4hmg
eRP144DS+6WoQ7Gy4mNE9FrzEvIX9L83copuZ41mg7GvRhgY8gN+kTqPyLo/PAuWt2m0D3RI9noG
kOYlIB0ccE9jgRnUMmhuLI539rHwjoAVuhBVeJpvhx+zZ45FJ8XPVX09nZGl9G+PlQv7oaPyVUOn
2mrGfa8vw/C3Ro+SP0V/W7+5q4n0UkwIIWxiSoMCIJiiaoyTyySGn6/aeacJVsI3UoesuEwPbUZB
WCLNoU/UobSOzgm9KJM3j7elJ3UDTdBBiCJD8+iYu6FqkjBoEA3tzAGzspOvKfWz3/jVkCIZkVUs
xfX1La77ZcvCqktsdxhFj8eAlA1403T9alzeq8S/Cvl+cQPXHtaLDQO120HGPEU1wSSj003/BxQS
UhuN2ASftbFpHNEVS5x7CJJQprebIfX2IiGofw5g5DmTe8mZIFRpFfSK3paK0J6xzTF8e+8DmxdL
SGTLiuMiAfRlu10488feHv/nBwHksVjc4NK1+LyCO5cuoiViQwo/K95eeDmVrVBHsGfHX9L4nk+G
TPnz2BGIeCo5R2cv+l3ZXHG9kKIQPGAwuY52uSURiMK6+2TVP1Zos2xLWodjIJpdBvzJ3k8RZcll
LTZln/+zhKhm2CTlqLOOnK7SgeAd+MPwd82kbVuVwioD99f+SUrqWpZC8GjILw+GzqZr2jQK9d1d
oAlSKu5xeTkFHLbsZXdzMt3uHDRsv78ax8GGG/R47+wgaU7cRg+nCy7RGcGr06iJDa9KA/qw6kRR
Yqn5XSm6DeYcvhkJGsLkAiFyverYl/gyA2rKQDbrxKrKTd0okSNcGbFnSdSV5xNWzO9aagVSIDjJ
kdvWwE0s3HZ6+KIx3UlrGHZABzZS+rJ6g9x0chpZLu2uajPLfAIRPMWIjv9jfWnP7ZyJsE+cQLHJ
guAuYl6xKKBDKUcj/Lxflk4Dg1T+uff1YRuD1Ehq77uhjV8Jtv0OetFWtvI+80xZzSpjBMBFGcZH
03Ov+aUHLxfBLlRJF8f3r/Ahnd8SemcwTme+IHXI1niotnK2+JFo+2p1izuPd6dxwgFdPGeV9vbk
c71CpBxc+7px89+Nojxr5701F83bI81bk5bPeScxHD8zQSkKbFrkdp0LQduSrX0m3LGGg8945fj4
+DgMqkZsu3OouDaHCiQvhON+APZp64/1GjEQEZZ7WewOzxGeQOUp+PXLEMq72WNNQvFwVZya8nzx
7TrpAKNbfEVC75VWLULm21HgMnUryzTOBkbRR9UkQIPYGbnumQTiOphMEsOBeNM3wwYNarS6Ci3n
wZBMenRxH6lOxKMXzh06niCfDToyA3YBjypOT+4KudjPphUa9JrLzEoFwoiRNkk8b7Vv7DYBFfpT
ztjxr/xULUZpf7yxa+eYxJ1OL7AOWkGDniQlDdq3tkVFQbFIvmg2oPV82ZyYGQQFssuLln9YPpBZ
Wxznw1ayGadHPwVqyVMFF1gyBwBwz+oPDTvPN45ump9jRai65+y/oV/9PE4I8ls09+TWqq1/sm5O
8nDLz4k7out1OXzMxPx0gkjTJ+SgtMLUNTtPWweJPBZAIudEeTV/QJ8N2x6y0wVvJ8MH00Q9uMUG
Clyh4W4j/lKzNELj0NRrcrHaArfVTKzB2hq63DNM1G605F7l65PqA1fjdJXuEQ2S6YRC1lSJ6Q5M
hA9F0lDmMAmNqtzO4wF7FcpfZiOkItO94sllCQN3Zw5sz4vbL/G4RAdkEg07uFUWtsgplkTQ49j7
r4QziFwZfo0GV0HSJOIloSdTnkJaVxWtBiVl2UjBH05QKRqKhWr7wAKmbTzlouwo6vmCSMjq+qpu
1asOZ8HXn16wGzbJIWNEuuitD04nIg6h7oTp3hjICXTdQC/PHuubYlrTBnW/I/RMlrE6UlujKg4W
tmxnVzguX2ecCEEz4H9t5qHbapdqWsLb+D+VwltjaTXukC8L6qY1xg896cBlHwq15/2sh1DVGcDA
hgfA/QQyqmtGZAXvQQn29CQVJLEhoJw9IwvUuveYhWIq97MMKNNRDDN4fXy3B3naX52Nayl+q/nz
uK68Su5IteofBuV2qgLdx9cS/zACXdbpyoj22QIkg4F6043TWas+Tz7CgjClmJ2yU9gpY/oauFFG
Yys0VbAewh4l5Q8MLnCjsM4lPNmHS7Ymn0DdIOGcJxb0SW1BLiHZbLCkPe32GxbdOnJkpeiQ/uaJ
lFPyueHIAF1FKcimOCrvL/jXjbtDC/qz6rv+WWKpniQ8th7gWkMrSBNCO/+8O+8IWHGm/553y6Ot
ddEYVoDSzQGtxm7Cb1hk6UvuWfHRLSmfvgsJDCg+T2JZzV/+A+xg8XVnJwIHVpkb/ROeOOcaT4xj
5Hae11ATVB1WAlgi2Yv4dDtzoijLJ3yw/3/FXPiRsf5W3bdNltcRK1acOP2grJGvIr+eW+zLOhsL
lfhtjXxutTub7mZwyQ88LVOiZkH0A1SFiMBA/K4c0HnuFe8yDkv366ayEac8oP2vFbuZhR0quMiH
BRVRs2HPo21iV/N0y6YFPbuaCkwnj8rjSUn/iA7uoLB/xMQd1h846Qm70h3eC5iI5zaw1rX5tklq
ei6G6bLYKKBeIzokE3FMJiLdYpZoHSbAJZBoIDDic77STnKpNElSivwjExv2nppg/vfGz8Tw9gfH
NEBnd7L5I3zyhzHbrl5SgJyFU0f1YTQNZJlOdzAf5UdfCdDx0CVNc8wjIw3u71LVk9zphdroI08m
yRL42rISZkR89cqkfuwua3PBabYfKZorgJOxnShxBQnVctp2hn8WMWONkELmwDP6WEUrShVcwEZI
vePbYi7h30gfwhdIdpYSJ1YRHjEo5pk42x+Xu78B4qDOxCkGI1PeVCNzw2GHi4eWRVEOBhIUGuZR
qoCmdgff/okM9FDpU7oV41uGdSUidi4+W63S1XxuSztEXr2Eyco4WdIqFQkL6ExcnAu8qpg2tBM8
SLc0UL7S736D10OqvrXG7Xqpcf6wpQdBI8RgX6kgHemyk/kZ4tLIp6vjqzGi6VUKoiz1dT0BxCER
0t3E3d4fzl+YjvP7dbV66YuOhDRDAxCAoWdkuWGy0MaoYomR+1VgMbVPjiBnWzKxX2MXGKJefhaF
6gXTjQJNXqEXXt1sJ6mODZ4yP32sHA1yT+EdxiN7HXGdIcOhFHaWM7lrGT3b7gzZh6hzoIWGyOgT
NwWICO+o2fkY3tTm9l6Hsnj5mxbcYb1r/cFoPN0HLjt1pCy7eZEzWZ+QAKNq/u2TnhhmaiF9YShO
ErkPGZWQjSK4OcdOtAoGWqZHLXLO4S92DSKJOFFSNS/WkDNOeXc26nwb/NJIWK/OfSdFrSFK20/8
Z5gD3pY3W7tRXSvAduFef/sutNsNF9JJMCx6YYA2RPqjjTFnfwkokyIhDw6fQvhBmF1nERK/7/4Z
NkznbHrhQotLmfx7fsWiVQVU2nFje+hjKOboJCjcsxozHX68NU4jph3HF2p/uZwby5DIjthfzqRA
yD42RVJRE7uw84/fV82kUc/TsPfKzgzEkJwc0ipY8ljyB0rZL3ziWlGJPUenBFgV9anLM+6cdxaz
o7repN0H51dyJ6AUlV1j57Qw1NS0qh6qp6pEaYomiQsux1epCiyr1ptH9QnBniUEgOJqJteSKj7Q
bx8tvEaGVnkLzYnjCJVGv3H5+GUdYnPJfCml+qe1QwvbAHLDp3ZCnfJaZEnqw/aWLXruK9poNpZL
nda55PNV008L21l42SpDbJsS0MExniw/8DANe7Vi1/wjPvh5Xpd0OwYlWcEF7Z2v16i3FfNy0k/v
Cl/rXQQb4fC3bHO3ugNN924CIH5PLyP+rcefF65up5OQHCSeWDlcMkrLN/TxwoXlWCT84LbKb6zq
AFkBdlgZ6WPRh8/jCR80LPlHyvhYxheR+uKT9cglKTs9t56BGAxTPex0l0Vp5tSRCLQDgXKBS9UP
5gec2g7kFd9LbkRCEpieEy+CScLrbhh4sv/lr58XXCSa6e17jFiVDfaq68h+unRKiN3IlJajrMeC
yDkd6L5XinWZiluKwvl195yVepX+JMnMIYO/kijO1x9DBkFqrWOeV+vUokKttO72nhpgYBOlyJLp
xQW2PDR8mq7wfTix+Sed1s6Pl12u1zhxZ0blcrlG3KefSnrtvnKqMY9MXxewxnTzF4d/VAFU5gwD
vSEjPknBV8muEq6cZt6hJtBLqvMGPvlN8mcd6bEZyuoTn1TFnm1Z+xoLQ9QJnvxdCo1233nxEXGA
G7Hbtb4biAaEgy6mJG56jDlxL9kLvv1HTCyN1ZPdomX4e4tqQ+RtbK/qJaE44RW8R3ZlTZeEOEc9
otxftcfgC8Mu+zVtRQ25ICdWomssDnm/pIWfaRxG0diUn7efd6aRxB2RiAVe1dNB/I4otBMXbHbv
pIAURlP3sPCCwNXYbJVoeWTmu60BFa+TUR7J0xlf85lBFGZ1ZRfdMc5jVKXXL/+oZnFdg298MV2s
Ni4zQZan6kr9RCf3pVu3e1xm7XOl9kIZZzY0ExwYqSawlm24HCMerUMLD08++7euIbLZdCNjkRr9
nlYm9iVxTX3L5HxTZFx6Ug9l5A5y7RjH+6/JxX/Ccm61rNUNYhnqXH0SlziU1SGOccWdFf+R6IQx
AHC4nfbZfy8O/CTkNfcslIC3bjEWNGmSZczB7CjsjBqIJ5pfyjtXAy87Wwws7bpFRjgsi8A+xxwC
RCFXUjEzWr8vopNhhtIA7oKuX3neXFmbCqPGk/5T/OWbD0hkwyMVRBZrdlb7r7haS693fw7Ab2Gs
H+DkwQtpeuuEf0feW1yXt6epypqr1S8Ds7Xk4fkOm6q1MhrQERNEoWsDEpAyQuTuUM9yw/1t4Yk2
sroMWhcE/SbfQAWndIpCcu9gPnO841/sRYowvzrgPPeGZ0WQer1tHWyZP6yUU3aI2NbAx5YtGNGv
f7sOCE+6r0o0oF6Hurht6GCDZpPnSoN1HzeVFAZ1u/2qZGys8MD9r+vIqC2wOf4rhvwsUf9+YY1U
BI5/nrJwgX/stCPG8BspUevcst6CeiTiWeQL9vQlIuIZUEQBa3MvBqMjsl2ZoLHpKDT1gBoHNUAw
bjo6kIGbCtEOl4eribDwQ/hiVJiL1/EZlJmCztp3ij4JenCk1/gbjyrdQSbVfnRVzFum5jqW5fep
fwErIOacV5NRTxBCZy198e9OqdXApodRAnA8hlVO6eiGJyQwEmac2ZD+Qh0KuHDtVTyUk5C20Uo4
cCIGDreIpMDPwY3kghO/wgXB4i/xm3KmAZy0slP0qzocL8tbbgQQL2PqQtkVDnVob7Fzo+0VYlc3
dshcCxvK2pa27yLNX5MKvN068gB+Oe6+CToHCsqh5H886U2NjQ/EupcYbEx7K1c0cBcRA0mye5kn
nwPhV0ecxerKHdKi5c53t3KTc8jRmT9lyDA2H6ajCi7k6phMKBLa4Zpg2UBKz8YfoLHCmZtlffRj
MnyVVLlQhZaFYcudlnYa5GeM5tzvtd7C8tVJVs33muCmyekFJCbs2dbb9X2hP16rFBqDPz5M5fhm
7k/Z38v8urMtsZqVmiWoyG5IBuJJh4Ghk8qtRNArW7P+0i/Ig+ujAWn4q5cTFkk2cUhx/5ljhyeT
VQr0Km1+E5BNpSIjbo/QiMx7W3qVT5C3C0Q+eq9g/GVo4hW//JQeW/eDsHpi5t7EivGQXQLGFhQP
Vxddp79fv3XRXqSLRoFXNvU07imjq3pS5twyHhoU1kPp6Huv13WU2g1l9whsOk32CwQL+4zQqXs7
JkEUuO0+ZMhletuo85zjySi9MNlUv+tSh6Jghrw37p5NdmnyryN0EJl5qowwuYw+CheBWsNwj83D
Hz64FQ7dQtBV6HcZsQJ2lnTjhXMXFNgxNJ1vHJWYYzKU1YvWxV/K/Tb/3RH70O4pqHK+jnnX5pBo
e7WTtvVFQ/JygK+jEUAJ8XYoxOoic81xlS8yzXMAKgLUbKwJPq7mnnL6oNKD/qQWD1Z4XfkOUfBz
x2kQrz2tOZYsVH/CPHwSbuW49j/4tOguNjY+WHsqtx4x5f88HNanf0ywzcdNAPHd2jEC+DPcqlpX
fQF9ytWXTbl70THmknKFt87piZB5ynBEssMGG49ap20+A79i5JlsWkaV2GQShKNe5PGK9vqPYxKY
QUpZXZjBrZJfYDaOjPziHZOkDuHexnz2Pg1MpXvFB78l0ZuLiAJkSa3XkIUHOtA1UlF7UGJk/+uk
Eo5AmwG7GKRE9M5yv7CYPgxz2Rlocitu56VJnmiYCnfHwA9ThFacKk6bS6fF+auEIIlQaa6tNpMa
zBIvU/4OKUeEx/Ou/E10BBEfMlL0PPjeZS4K5a2WBE5/bUEBBW7ESwivz4JX8fQp6E3vhc66F1FJ
ynkCeat1JsEirJ0KI0aIORU5z6R61ZxUmPffQ4aWk0mbJxWdZen6C6N8ZrCZb4pAzrN4In2qTutm
bWSuggAB4g5f7Ky3zSB41VJ180VgOp7oOhmbMZosABQFFUJDL/+2EjDICgoSoXV26NjbIgSKdiRE
IgNobgc38GHiItJmF7gpg8EIYEcFAv+eMBpTfK+lsi4GwBv46MeM1lSD/E89qwGsFtSy+QyvrBo9
7UZWv6xfYx4i3SZwwLwleA4fmA0Y3Vv2mpvNHUBrzVffUJ/cJFRIbrjGr4exd2zaS/ya2aLUc6Yl
h+j0QLzmPk5qaedFf1+1rbuZDPFiGd4i7RV5UiDbcrOeDsPQhXm4xQTy6UbqfDRGBSDgZl1RKzKi
p7hgI4XglaqElH8BMVDkQ2NoyAKl6AFD31voVmu31E+tRYaFlewUP4kPzOVnnb/4NYenqSf9GrIr
iH16dyfUC5nL959m7ThkRDN1lPi9kBwcihMkhoo9yjc+jfIc2J1tgbifbeRQU2nQkeqNtiByR2PS
tg1Upf/U8JPcahwligxcOaI9qG21cyr/7kCnPxuKH+RVUaTKeLQjWq/kscELK3Yjf7rAOpDC6hZ9
iN86b2YX/F2B7RfNlS6lcjtVEruPTgSLb1qSaHzAJq4/qVsxJaGut9DqyOhemcjIuBeKLontirYi
nEa8DkVawjr9VKGjWoCPoy79IaAGBe5tZkAWbdNvBHE1976C7RDYQemefX4Xg9QK9ffRWRhBfbc1
Fh8GjaV3rIL71+00oymfeTUqtk+ksHJaXJiS/iyeoc93fKvP4H88DLCiDN1dH3zdWUz4d7ZLdYcR
H6EcPzF2NLBy83d2gkfImZjjrZuqlD0YwpiEdDCYoB3E5TRFgQ+lZHaDFnVtMgy85mOKWfDg+5y4
LvmbsvzyPmYxkKyoSOkvV6mad2amBVUU1v0NGN1VawcLe4rZz6FZkbvYInpU/tylYQFepl+EAXe8
VjvSDotQEcel/rfvGHfnWyJm1i5/CDVVSgw5598yZrE5wIQ/haGlM8vBxNyitnK8uVCoAuvX4sCI
IT8Rj/AZMQSgwf8udDn5TMeROloaM6tpncRfDKjc5ycB+vsk7RGGQSc4DzVT923oJLoSufI/Ovmz
bOH7vTuDZKzSl1NEpz0aG+xxhkmjRQtaan49Xm8D8hw06qnKP+KN2L2lqAQC+n8kLL3KI52kbjUM
M+DPiIqEQbteweJrhAazwQvjq5TXnzMUff49z+EHRv1cW4WDUqe0vz7gUfTamhPMABkdtSnrJjll
ZToOAA7Vmm4sVNfFRhSgxQikdNiY789uo1RQ8uejqUVu7YBvvbeSHIdIvMpbby+bl67v5eNShwXW
JyW7yGc2tJ8BNTUcMOTBxczPUueVoit6TtnFNvMiAuGO5J44QEAtLKPkw0j7u59O1OLG2IKnah+h
fk9WmVT2fcWU5wSJRzEfCwYNSwpO1/2fk7AYVYQMGAQWMe5r6UEbE6T0xUFnAI86mzHk7Df67mJk
5E4qEWbecNuCHYZ+NKBCGbn531Xf3mf9zvOHXi0JJWkdsrselQvEILbJ2GOBZqJVt7QIsfjuVkOG
oDCAMkbCD0NnIwB+9HuOYy/Hjs0UwrKQNWkTBaDW3Lu6mouKofkaJZmkhuemPTnlnZdnIdTSvwm7
BZSOpvVDEGyABkxkBxN7BofBA1iPA2RByRY0pXFD61kgmnXxBYxZ1CyL1DWkllM7+KbZ11eWh4NJ
RTv0nwD+r0bMjrhlYRcm4x58FP6vsTrNeE/rzc1MTa87MPkZrQC7YMDBwUw/UvTNCMMAPPjPmgH0
4OdUtPVih9i6yeYa45qxPXO65Ik/AR73M1/goP5Rpm90TMoSd0PWoxEpXpmsA7gyd+VliSRIxIis
egkRsdWobbFKOoBYGcMRPcoHK85JCeagGx2rdRVeqP/jegWTG64DBdZFwF6urFjYN43BGTjIR4Nh
KhxnsLq//HXg7zVMK7LMYe/qeiA1TmtRwDTc/RERjE2m8ngySLL+eyTdcNfs8uMLpi0hIw0dJ/1M
zQbwrao3R2ucCVJI6ufUpCVZMQGtshDFCugI3Tp/4liurgmOn3Qz4j24sEtvQPXiI22rHhzn/p0L
PKlsLXkZLwVqOEFnKwgPqJzE6tkYrxCUYHzBQaCbVljQRlBNLKhGPgTA42F1z48SeDGrC0gTCezN
Q31Mjf2+IenjE9amMVBfwvCG720ElbD3pHQu3MG9tak4WB0Ps+p+zg6md5qGHx+RJ22Fb9+wPnSo
GRmnmVRfWwE0s5EnHIM4J1QpTY4nxVIFpDyFuvUKA4lYfuGD5t7Lq4pgbOeXCik6RBFvXIVe7OYZ
4enW4VPP4kCZTHFN8NHDsOFr/Cg+NEYsjdO4XE8tg+JT6kmj9Mz0in1z+GJo68POyLaGVMIoIRxL
kD3T4HaYCS7AqlYoWos5vLLXbCn5NrIxjosvGf4BNOgsoordPlJdw9qrYYVkb+DCwUkYLtQtgyzq
9cSYYVvly8brhqzBsfWLpSmaXnx1+zr8VKTz8BSROY4/9C6lATKE3dfX4OfIVOzdUO6iNh6+L21s
0g2Plcwm27tEXL5FL5IhH60E/H0ewuu6YwBbMYbxrces0CNfNYXnNaz1C6u55NNItaeKTSTS1sBM
J69qlIOVfx0ie5h5TPgsfyL2lnKBZWwZjkvPZQJMBUN+hmwjEXDx/PnVEXvGLSRzEpZwUWd8JHSz
2GODcaQdJ3AJyt/Dfy6ViL/QRtqCS8+jBMoBlSLMuBeaHLx9vs6GToagXWTM2h3z2B3erFeP9vQM
UuvQIVYB7fPM7VghgEHNH48Lp71uyLzMmOT3K1fY7rdInO/XinbL5BUEQV4yk+u6fPpweZYp7xZU
PruTFVY0Ir36xrrV+Ks71Y8dolgY8Vf8DUH/O2aUMykc/ARHcXH1I4sbj80+hWaKSjqBEGQOR2eI
zJGAL1NhYLFB7X+Q68q4lu4FQCg0W+wAkM2Zp1sBlyvMWeTHV8eJZvkPMz9+Q8sjp7K/dRaMdONE
/zqb+NvRrL8eqSWX9mPlpL88n/ujcrzo44NXYyD17z6h4v48bJVhmHIN9k7fy8a+rldSRdwnVHXU
7dZ6pQD3abRQkfwcRyBT4DlSZfTh5hnTL+FBSyYbY1R8DcgXym4rzIU7RMH1Tstjb8rlzJLcNWjt
GNHTHCtm0kPWDZSjSbKcFa0pTc4Wuni+9X6/bbEExEeC5ZGsWY3ckB7p6eqrM1WnWCyFGKewAaFn
XwrTb4pmSaN4CYa+qXgxJb09KE7RIk4ug50yFIKibRI5/pEv14pWGLpangN/Dp+s31kpaxayLtcy
7Q19sS8hYCrR/mc31omEW5EEoO3RfQFpHIDttMGIxCqc1dpg4dtVIHqRqV+HlraKaERn9NezEE0x
hFe7JXkEEP/XE1Lvo69c1wPwDCmKAYSUBip00dQzUQorYmp93VPlgOPb19dzHLH2G/c9mBlL8pZc
p4xntG3bL3OKQiSqJJqeTswpZHuAqdw+YJEXxiOLVnmFI4IyIZU3EAC1x24fyzkTd2e2dYSM3F3N
w+o2NSrehkh3PdTKbQhKQ+Eb3PDeoQ/zZVtUWb2Xf9uOn/vPqTMf9jraEWIKZlyE8JK7z6GhWIPH
sZlg6XsXQmpkflLjH1f8mtcUwL44+HoXWr9DhFBdVseHJ2IFeiuFjfTnQwWXHXnII3UBxQMG/JCB
hu4cJT0Pnioq24JJUAX3uKHyc3Ekrlh5MP4eCMK/gKLbvqZpZTK3TtEVy7FEXLqTdyfrIoJQK0Hc
XWphxKUHaou+NWdwW1XpzAKQTW2bsWWkMDpbsZbzG8OaDcoi/AGvsDfwwL0D6EpmjTfB4FN4xdk3
HtrKv0YSiYMKLrQ7k8vLSDMHW9XCrgTIAYRivISWj5VomnzNg3/H8NivNaxyB+r8V1zuPjLiN/Rf
h3nNtVh8Vxm2Pua+L7o8czczCV34eRIWLbyOtUGgIWwZ13xeerz3K7SxVJsO5zQCAFU3LH8MFwEa
mVxhZKxQ5OYkuK9RSnvcx9EP+3cQUnnEKgYrAirG9uhLPJsWOg6H5M5nlL9YuhHAtMR6j0+8Bjr1
PuAowC+K8JvM/dnfY5lrydvPpt+/rxg5xkWk5rwWWl0GoM1R09eQ/ibvQiacsdUM39ky7XCE6+fX
ADoRKFjS7KvMH6n15OGpEy7eJTE1HPIFXcZYt0sIMxu5pyete80hHUY7SPYEbJ5nQktNOuQ+feF4
wuy2MbaGnWHyoYzMfBGWBtXpJzRiwqfP/LkYjB6Z91l4OiI5DDAllDc6DrZj7RQFTytA25gw1otP
84XtQQ2CWWz3b7j0ulW9DYDfkToo7eCTTC8KlO5E0iOdC3tHB7eyTx4TdukxToPLsexPF6LIdG6p
bjqd37481NWeIPpDRn8YbbzdaGzC64eH0yCfrQjjBmCQkqe7JRexSNzLq6u8JwvK7WMCwzOneIjM
n56Vk+oNtDEQwboAPgnjyAVddL65udcVeiyCysen7IZBXgvtuIT51tQzKhQJsgG5keXJ+n6tD9GX
pxSvJbR8TDE+Ah1yOH7E0zLdmuvVBMhPDyqlExXGcawchlw7obUUr1i0K3ZR49NwJaGHLCIF40AR
g05dxzM42C700TysRtazv182Cic80+idvmN91AyN4e4cOS/lOVwh1xJn+UR01ZBsoSNOmG3Cu//t
UtRgbQYr3cgkiNv7lksGls2qbVavBHXYXgxZyLs3BUNTcwNrIx4ZAYEXUQwUBxgkI4mOqC5rb0nh
POkk9tvH32MeKHs1Yy5zQWzJ8D/iiZpiElHgaDlKU9ljNHX7BCiAH5PulU5Tl1n122LgXvNlmGUb
JCFU1iqyAzdNxZH15LFxMMxciHQaxJkhTbvbF410ryVNAm04MMuT/8sel4cS3J6Mz/bWJJXTjMV5
/aqSeR6yTMw+3UqJy3HhYoj95R44RhFJWhbzNB4gBjO/vf6KtSNJjbBzX5+9jpgVOumaJV/Sf469
MV8SPa3oU4pafutarEGz0SFUGGUINDWgDQJdGfpJFIbsNaSPbP+ypoi9i0FGGB5yH3otEuPJwZ8Z
qxlADTZiSb542X8DIo/Vcbvt6tKzNoGWyIhg6eJSYIvCCQ7qKu19kL/QjIwnLlNsKQqhGypticmz
9hwnBF1BuieYApv3+411s8V2I+vCWodB7GVrJnLyFu29ORL5WGFX1aQVE2s3LRGEu0fwenGJiFfl
+jE/wRf4HmcsQ932EUPRC4lc8h2Ic/Xi/OZflET1pwUz5hnMLRAvVydNztZj4tXvXRWSwh8Rl9Zx
zSiS2HWRQuNhlA3b1hHeQyEOLQhBQfytCDVnhkBe9tujg8wkepHXZ4g6EQUokV02rx7kq+Ie9btq
CIopRDO6VPbBEHyEmMxmIdD7+aq0W3ZWVU8qYouXbrt+JbsYvBe2eiYHlrJEZI9qH2feeXSivPMs
gliQeDs3R+Hur4cDoWzirZvyU5UgswBFVtqJ8UYj4MnQyVnC2KFGwYg5fP4KwJ45Shw5K4p++2ly
vcSdMqHA6yN+XKzyb8rKm5NoHBU+IZm9aXUK/Ux4DZ9iN0yUcsqpvnwLQ0KLZJIjds1xqqsTm5wf
B60eLZJMQPZ+9rfnaL+7ba8TwiVN3ehItTaoiHq/hcLkrLXw2JQ7onXcopj1yZdoQZ9RCuwjwRB1
Zzzq1N/YLqPajKYIYkNSJ2iU/beOsRHfkjemKDApXpxU+bxu/Em+UoNEvpOAaPFq4AnZe1PUa58R
gaagEfPFUTLaX3vvEVpZjcn+1A9GLXdgDHbzOAFP0A2xjNU6MVw+FSqWTqrsepJlshmkb9dvlUya
A8rVaNcC35kDs6uVFNymMyfjYCwOTREkSCbOM5fbyJfuhXCtpiGzfQEAiinHEii2PaxNnDJqA91D
/Sg9k64AMRrcJHN14S5l8ptUf7kIgnInX3983KinbZ1lb/8EDCHfn4UwzoVW6YLWnwTvRiyCC9j3
CJZGDTXyV+m4jYDiE1AnLBAl4/Auvl5Aq4xOKBA3lunFhbHe7fnu2S420Yy4ahibZaFEZ8HJaSwa
/jouBYvumHWjHHnrKNoKi9TEEgCMOrUc4Uwt/OZSmQCmiBY8SyJPlHGZ/WKxU/ciArgM3SYmPvue
TNrWYg5DmmeQOkT123+j64SYXyOnJ2QYkpH7MvLQR9NpD/IkpFxEWif5TEScZD7Zhf3XrTN3/XTz
YPtYijgqdqgERs5fy0zTUsMH/c6CZUEqVoy8PZW1ZJFj5nzt5BEXDfJDhgv9p2d56wAQmauQAO8g
e7vCT8KGL1PC29chQt4qfPR0WcvjYGAkpwj9hiG9dC11TV3H8Vw1zCKKX23eDXi1DCuoAGBMIafD
D8QGnMMY7IsD2a+weUri3Zv1TYlf2Jw4wduvynb9FWAg95fuezO4zJch8faHiU3V88rsJK5kWlCz
l++zK3kCRBiAxL7Op5Jyh6j0kdd5/5hTAOjYNwYwZK4eXbF5ohnW7jqfdQiWPPoRvRsHEQgX2BTz
0jpnDx5otscGbV/G9cRHzcWKDCL6nlgBDfVa8UISBJqcooi88WJcO2cOq0zB/y3qgeE5O4LYfMp4
Ivfz0CVflDyOjdnOKFaT5w51pLphNetnYCPEfcP4K/k0hZ20+KEFgKCrnGwwhLOLkIbDOlUPEICz
5NRH0YEEVGb7BhuCPn88PHAg+HCwsivpkPqp741CHEVGUqF7DJMmCi2UDm6VNEQC8CnS0wcSjdDi
KlCRMUCnxvtWEwZjqWRjoQoCSc/FFw3pluFhjG1azOQUxHoVsRhTgt8jOIgh9QQ4LSBh3L3HEVcu
G2I3jAKVGPdH859B4yLnMMsxAJQViptpu1p8bv4AvQ9+UE215ZLGeVrDBMVBnw/o1Xnyhw26YHrK
3RuenPyfm4bLzq+NNGOYBP1coFHovolLOketADMDKOhG3gv+34tu3fZtXqPCpKmqI1+iIb/xj0+3
IvfYGmMylQgYCtuzMShKXQ+nPsijygMdECf6I/ADiWVlVMtLs66PJzH22COWmSu+4cQ52WmbjJS9
/mf8xB9tiAWOcfc4cZMiWdMP3mrLFPSmQv2Pu9NiUp4AKinYsQwhvM2iP3vqI6Z2hOisUUUn3+V/
8E08uMV+9UX8FGDb/TLac72iY6v1Xh4qCYSnI+1R1yhvoT/WM918mNEj7BLoG7tErndrQaZtWgBF
s2nTuGnEVPItpBcmt2cDAMQWOEc+6JjAZYxaCqimxHyCn8wfqCNFR3MhFZu9qCWI6taX5GhOprjA
08KQK5JJzYj5wBiJaunwfK2vxfHyUZWzRKLJDloUHhFq0OGOjzNUb0SHN+D12x3mupY1KFWz+q2E
zRMPZ1XLD01Dv1V6X8dCWrwd+1BhjmzedO9PgLr+xYQDGLKt9j1M3WouZyRxgnpvCziuvb7B4duB
GZJTxAdyJuIni6ubocBdb7N52E+yNezkgzkvRKqgdB4+q8oo51D31X/7a9yb9V01a1tZcGZ6tAqO
ehmZOWei+22H34AuIKXB4pQD+Db9u5dDkj9/bjy4CWMVyG5Q6PbgcCZmnDnnzJWuf7wUksKI88SK
Pc3yesENzAgWbgd2sxe8r63B+J1Q5ONEUV8dtPUh1rwU7sfuFoJRt3yW9EddCO8P02EGZw+MkDfV
tJMnn/ueeS3CLnPltmYDSVEhM7uqkVlyiKN4QgcANej6ZA9hNDBeQB+91gzE1wFxlAW7G0891W1V
yPqxSaFE+cIW6gjT2u1W4IvQhYY9L+tEifoCP1RU2k0yNy49XgpZfk+OoI5rE7LnIsfBnBxzNeal
NgDLTt6ZQ8rqk07IpJT3eLLQSkoqIxpKP7oQG4wB/q+ayfDMojrc706I15xSawLw01Uikj0i8yWS
5FoKuhwSj/W4XEDUD1qnBTaPyjtfujiCEfpr4YCE1n997zm6TprBygfmiyZ0hdVtRNs8cdZDtNx0
Xquzg4O3S3YgsMFfEwXOLuLoCeX2hOPvbDmYJtGLMYtA/+IZRMF7XK+4UtF4A8uiQ0WoMGjtTEG7
M9MSwOfWoV8Acw2C/CsCeUkyhcUU+1XdjZejYHFgGNGp1otfjOHoE4tarse7Tjhvs8QV396lwbKa
wmGtDALovQiUjg9y4/oGTu9bIyzfvmSWTvVpxfFFCxdvpN8LZscYlydscyKa4P9ELHz7BAVdRDOF
p5eaOzbAFeENj+xFdqaUH5iMkbl2AcIGd4tmGECebfuJd35QiVmo/QTwTB2FbFtaQRAog9N5G0aT
oWJF6VEDUjxQT/WCGIdjumnHrADx23OcEkXWpQLR/jC0kLe5Vmdywke1qCl1OXkfuu48J7omPWZ2
AMU5C9zrRHXC6UG6c/Zecaz8o7RouiU51vv58+rJv00NPZnim/aXwgLg2b8oKz+aIOTTIWLI+Fth
N+31tMpRrS609ZeBmJTxt5fdP0mwCij9DZMbEUjNe00rohzfY9njXSzI9ZXySPGhnSbPo1yvtYFc
vefzYBQ+O+edyFl7bqoXNOmrXDMhaxG9pmIOgOG5RCXWMATyGWfcH7KfzNF2A49yyCqnY43rnHNm
tzrXG6KNiZCE2U/F+8T66j1johY6zfwoUsAtC1x1q1RZDCIaUaFBmFlXLgwuiHU2tuPSq5qlg5YD
HrxgEKm8S82yCuzvBIN93y5EbGIU/VrqVRcK97FkB/qqiG0lsrOaE3v75B3nogAQ8GY46MZn3ZNC
u0qXfVxnsaHdqFmcJ4i48cvKYvYIT6WRf2Hdhi5wECS7TdTxA7HGH44/Rvq1B4WtgAw3nVzF1y98
slhdTjqs0Zm3sWrtrzK3dmku+nkjq2A2OVC139oVWUwZgzRerXK9r4i4JFOelH9Jzq+T1Pj5tdDa
eMu6bHGUYesR/NtLAZAAhcou50I/9Dfgl5ZgG7WRFit5IProiSaAiU2VjcNxb6NanF/b3+/jsGJv
5OVi1aUR6LmpCMmoOYfUnMu8GvuzaPsASZWuhMd2AbXdM7EcvCoNYiq/UrkoAJPtRfJwRH//pA1q
98SGVcJAw5/deJ/imWhjeSpA6eazEDafUi7TJhkZ9inJwPjy3ByxFH3JSZrBSlqrUwqB0i2Xy6Gd
M9pNVAfqp0BmSpOM0MnwZRFgHfKopWq0QXfpp7U7tKl6U/KSP4Bf70dnhV2CUBeLRmv5X6+6Nqea
PjrU/D9iiEOPX2FPDNDcsD+tOaP8yRaDiK2frxq6H4zoPJWcj9UXfyIopK8PxjtLOpXuQP3oqdqQ
6FzRtYnnSX6Si8izTsOtwMFp5KB5Zxo14D7zr3UZyqDd4TPhQfIxWA4xSjZQ+FuTyNwSHCA1A9Hf
0nG4/AW2tV09S+P/fFbPja6s29xfbNdGBNg63k+hVn/eBVQGR6f/3ziKuULT4c7D1rRV0RxUej3g
zXCqYNfxFfUkRG47ubCz0QHP6fQnEvGS81LrfH6f/CqmRcf/dweoNa3uZWdKSrjJkrgp0Hu7/giz
k25LfTAhWE5iAyWlvbPQVVbVoQfbmb5jXneVinFvBw8WNSqGGVVaKgky62Ws5Gtuor/8Z0JvdS4n
e6/mxmYibKyL8ges0JxCcj3fMLJ1oysF6qN2GpisxORzP+qaJdyGbX4TwJbXgcjnMDKM1kBc42z2
FAPQJtoA1eK+vKPTb9QL9TYd1bunXJa+HXSnD+Tebs4DXEToVN21ZjWYiTSGk1CiKW4woNpPMITd
BSQRlvi4SnwvA6ND/Ir+qGkAq6vgSev1akZ1QHKjJ4DqIA9bR+1vPWhViA0DGeIhosoBj6yZJA8z
nyhk9Yl9r8oU5Ki+mWzN49iRZ3XPtP8v95zV5R3hsF1pxDVflPXuH8Gcl2je2OAYTuvnaIedoGz4
zNBN/PpWS9r1RAbSSimUxgRP5PRKrzhDejJ5BLcRglKKo94BMdobUgvywiHaTUKNrw5Vu91FueOk
QNFrzO8GWGSuImjIdoME2cM28O/xCKQMUlpkC8Xq+dDxby3QYic/GrFK+2lvUaU8SqyzMb8wlFOZ
K6wDMPzebEKQHxEZf3BSchiow33GAyjSV/Sth59Utdlb68pFzdPk51600YF6UGSvjjSVLSwmjwoM
d3bsDkD0I9U63E/1LS9gJmSWr0Ktc+sCYe89hoXbKT4Se5RCXVLVkIn0aQsB0ak1zsm081iL6tnN
qY8OSn4drM0YweTqYZehMeZffDHBOVmdbstlFZxKocDqOcdTHGMNZJL9dFs36rdSCEesSW8uZwsE
L8fFjXNwhj0GGTvIYyDTUBBYabx+SUTgSTF9SauHGHCgtXZFzNPVgNp/bKxbdFW9qt3qTuXgrQ0F
dHmXtAsLfF3MvC2yCSP1TERnM1k8owgDrKOJIrh99PyUY4MzRsem36mJurIA68ElZ8v54P9cE4TU
m5QOa7IL/4ZWhxTHDwhZLPnuqYJBnTKiIiiv28uFfp2wEE8OpcgxOXOtgUPy+IfvKECJoYN3zGYq
A92kJ6SoM8PhXU/KuWzllOtLOqQwos7y1FA92ER/C9vF8De/2edLw626FPpqPDyXdoBUccNHmgyj
K2BPlFl69wb5oqC09DYC98gva0uZINhMt6Uad5nqelm/aksMVyVRgCmurZLKUxpf8g/vl/7DtZzX
2ulcGO244T/gDXuo8x3XWOi2boMzjNiMMMkYBdSJpR0b67+sL1bTxRnZ4x6ZOYAZmeIU5dDE1L/Z
L32CUHGzaduVUq549v9M9qsYzk5PPDs+mcJfsGrnBYcCsaz1CCHjlNJhZ+2HN7LpIUCqlxB/UtJC
V5u0OfRaZN5wprKg4vU/pQCXBbm/EiqAa522sUYlyt5w1n6NWf2YuyyUBDQ7IMnuGSn+Yv0nIW9b
HJJTQpF7kl2VGNyws4TmNkAVf1vwhHHdIxfYgfM/bKGeZ2UL+T0cvbaJ35KKyrlW2OUxjlavQ9n6
HhTUK49KDlEjh8qUW9UUb0vXVqQGnCF8jt/Pbc5NsCJ/t6ks5G5G/4bWaX0pMWtU1YhtNTCA2FYf
xDl6BeqCS6HcbiNiAaN+44Nh3eR7+FvxzYgTTYvZY6NlH22fB09F+nvNGx3lmSt6m+OUyFi9rBED
Tqo4MKexyBXGma3VovMZWjmvOhOtXgMYYNMJZjlsns+FrFW6khOm3Q+igMlv0CdaSOtTL35t8Mqf
FnQRTxYFtoXA+FTL7uoK12pE8GBVT+0/fp4+UwQFG5X7cClxZAVWZf3lNtTC6YboJdG4P60zRcqM
hpWPywhdA+H2yxJCWTNLKcAXEjSJWUn4o9v4RMBL9zFB1CE+7+KzZqMGdFVrgVXsGXnom82yakMO
19I3B0hj6mJFiwQzRxCcuv/8M9jv1EWVhOvS0wJGUEbfe1PltESZbwXx+vQhIYaHnOA+qJ1U+PCs
CZ8QTyY1YVEh9AQTKrvpsSi0sqDr1teajiZm1Fs2hBhziecpsFpAQrkztZDOPxrjw1+ynLGv4qGk
Mp5NN0RaPoogquxa83cG+uDOoHFdUC9cGbd/WE3pRzoQp5l9Bje7DQVO/PYn5evXdvMAAIIjbQwR
+SndhMzM+BCLM3Wi9wHIhF0Ez9LwLVeOf7MP9Gn2vTfYj6zwLd7oVaMqvj3GLfoWqxZlXbmG9lmp
dAHd/d0+4QMOBOUSL2jKcbwmooVvCTCZPGBMbX93Y5VpOmC2XwhWTXqHh3oxcVObZc+1Qy7cRPbh
aY3TrAf1SgqDmQbRn7KwWWaemh9IelvLM4JuTdLL9DZSSo5r6ad68yG8AkATYQjZBOz0sJMT7mi/
doQ386BOeCtMx5IBrh67EPzyBqi1AHcQN1PrhEhk09v36H/yc4jmOiGulDTxJWrtjXeRX4qRVh7F
2cV1CxtOLT1ElPbpHiLkGO4nDBK1rFNAHyQBY5jAT0CFzFo1yp54XFRxaw4yZOMprEL1RNAjhdBp
rTMu7AGDQFyzipJa8nYixG6ef4+fBVBDqQcm0IPPy/3ebhlw+ko8mD994vO45u8Q5wcfBY/Pv2hK
5PyeE1gk06Cig3mwKi61Q+seBvU59HSMGG2c+W18VHdjlZikS3TfUcLZoMbhnSzcI7W/IN9xcECu
2QNmmDeBA6uk43s2j8aB1a2jbCRQluZkaZq9kTftN5tOK2d5qhQ+dK7XznMAqbwZCnnOJde+nJrF
/SsGyqfukvkOCydJPqJDAg3ZaEJuTwkteHNMOrlgs6P/vRBtfwGgkwbVYnlxi6tVfMAy0pniRSFi
cZ+Yjz6wqr0X8t6RKFPbCJUYcCzuG9jv6jFHG9rdeKPVM4DE9FedHoGbj/Y2NmB2Ff3bN1KJ1mGV
4B7mrDoLeLcH7MeWJ7l2E23gnTN1qtj5/Fk34yLes+19p9Pmhz6gCQA+3oEgIEMJL7P8tKLbxoGq
qbb9OLp3D38AY0A5eap2H+F52iuxaZVbuRb5u6v75QGyZNPIvJUxLu8us2UcKywLF2IWHC27al+B
z/lr4biDXSIgyv7T8k1zMIsscGEB8d+u3hTM/qzW/pBzoVibRi5CTHEiJta+WZTYG7EH+kAXwiYW
o7pcS36DVkJ8kF0QaJV4KO+/vF6FVAjpqJ4jHxgftoTK6eET+JLmYQyiV2VGyroWj5qu3IqlS3DT
sygLwTH7EJyg4+J9uNqB7Pls7KTs/CMtYD7t8lRYgb/jSuhKjmmFUFOiZlAIFyL3U39yq7Dw7SFm
S3bpC3oxU08KmiZY4MBUBsvU927P5UoiR0mSIAovyML0vClBu+h9rK9E0Z5N+Zjbn/rcQLNQkciZ
0M4N+CJMd4SxtrkI+xvF9eYCLAAaljtWN49ql3pyqh/b+mGAw6XAjePBREgSUjRlKZDpoMp9KEqy
dW5z3e8d4maAhsjeDjj5rBQDkS577py/gH+CRLhdp/XhAGS3wuz1BlJaAsA4tnPueKb3ek05l9is
tExLRCYBWrNhxsS3yLmSqm/uAuB0/aG/9LKqYIkogzNF93kUBEIiGAsjbYh+qh8bOdVnlQNunPX2
xOX3TAdw6iWLjyqfXp+BoXNpFtUQac/DB5l9xjPXbYvyrgQPYb3NrGAMM0Keb1eFdGWaBU8V3On4
8s8hSWxTm2uLlXeK7QS2mIWm8bPS8+fd4U3dFkbXTVwpWqQfLnlrdxqaBT7eu+I+HgkhnWH6DtIE
B78vpWiVtVqF/8gbIMkllS7BE7OvH0p8OD81/1va2RA4QUxRxmTafF2AP1SFm+P12nCJnekU6xa3
rZDCntJFOn0mQZubGkuyfLfGlMUjouXoVWMsqYpolWs5xbIkk7/2b7vEI6rU4Z9i0rS6aOf3lydS
+3CFPVSrvWoSK6+OCwAyxYtXXmow0U+gB/MC8/4rSmirDx91j/J3RW5SxqjUNdhAriGDV5uqINLK
a84qfOPAyiR2wf/nVasfPf0P+J8qGPgapfbY6P2O+rV/XD3cKOOpdJyj1wzFSRiburo1MSCHWWlx
nXlTZNtHuHka/E89bxBujNU0ckkuB0CIJePnr37glPv0Jz1VO57W37H8V0yKvEU5Tzk71evWlZ1n
tCCZm9PkSzTH1ckNkh+iB/gDE7xIOsJT8ymv4g8Sefzio3rB2cQVGJqtOMz5Ob1jMuWNPDg5EJ/9
J5z7rh/qLLEyhZzLAGMCGyR5BZoM7tJpHE+dJ++xOALnJPZzIGNZLKWbzdJ607sqvXUbyLzyvJU1
PYoSXIu5CTbeyHo3HkQGcDJkc5gSZIwjest9TDoLLSRGbzNvE5xcA2iyYGlQHXZy8TS2zVVqBeR7
jpQ5OccwPyCO/FyQVwMrIJlaahEFC5Z94RBw5G9MkiK9suABExo9xZHBT1tVAs26IOsWdgUUDIZj
9hHO9TWN2w8YPo1n/hE0gsSwvnttWvUwtMMEx9sl8y0flBzVPschz+X5vFXckr1fSJ1Oxaqv4vTG
u69QiV/vVr9EObESfVZLOCxcr0DQaIgcpNFvBLhTZAjIcU1lqYMrNq4PHDqwGnzNLUX6K8u+8TAl
kKfhUzj0nS5+6Tjx90xXv9kDKPFSpDuMTtbh4Kk7qlj0i6zrH/srKxkLuvv9gbxmmHhp7QMUd3Ls
s48s5RhKQYp0AsYQmyDKqtacecFaqmlNNZJyAJ1ra2KhV9mJTw8X/bIJ5T0+MkYWbtXN5qsrmM5w
svQwFryIQrdLa2bj+mrmmSIPoxh/RTbXcqhJxJ0D2SkAEyOqa2LXVuiI9dTaHB2zBasRencAL0fc
XikOTv48qTZQfQIqwwhmOCOmlvL2NY1/SylF1e4A4O3Ws1Pqt8iyHUel2XPYHKIK2tmSPwbBU8Z6
HYpQNPe+gPXKRAz9HDvVRrtdLmMeVyBUMUa4xwqrzspZ7liHypLWtO997Q0ulxRMQiNA8PYmda6j
bRlMfVz0Sb1RGEnCyLUFk3nEIX/qtsTmnD0hfMsH402HrBF+IyFBdBp0A8rQWX7eok+W/kmRmd7P
PPQUHxXL/gXm14TE0bdVFCOKSEFcPoP0d4XgI+M4r8xq+gFrFvUdO71Jy5KhyNSMdPJhKmHk+P/G
wWEYDH6kKOg0w9pDHK1zNQb7mbMpsbQnlVAPJkogpUgojA2ytvL9pCiQ2i+87oe16x+m7Z2uhrAL
aLaeGlWMLVkjD3zwj3ayTn2fajrk3qwIZ5MFavwZcrBNupuDUsQ0Jj1fud9a+RVPpMe+H4Oibh+9
UmpWN/zJtLH15Emygs/LipDIzOmpzdMuo7qK16haevGOfHfAtItPRF+SXlCsYkYTOa5bWQ/dR0Rx
sAaNXapYvCdtHHERSsN94gNDCQfz87Jo1tHpBgY6s5gChKC2+E17MaCeoPpovFocTBAWtOlZPJI8
TjEhi6xFQ+9KItBWB6s04MkW0k4hEevTTrFhE9YtDXKiRzTXA4PEUi4ng4keWN6avKVDcHvlY6qg
GBvkz8Wjosq+qssOAZDxfWtSJccuYnS/dABMSm/wMiiYLl9ixdFAhE4mTrLuUpqyw9LmDmtC3laZ
MQmsGlY/iJ6GygQ61htUzM4GkkxQAyq1VV1W8TQEv2kmbXkyo17ScSbjrKdN0pza/PNe98Fanrnp
zOy101xtE+HAKdV5jq4wjDGVI3fwXPHq4eU6uMXxX+c4ZGpVTCKE+cL0/n7JnlPresMCy19cEoqb
OetyUrbRs0ige4O9V1zfUIP4/rdjeczxD96D6WEljz6HDLXJgFIGY41MCzZlGC6FHqgd6r0vYSAm
PGHI/xE667/CI+NI540z+OnFSME4AVSW43VZE5aT9AoIMlXn2tLVQjK+rOGlFe/1ipN0gKAt4Wr3
uOIzjOEZHtztJuKIAFPs4JszsEpc+uDT7QgRs2dFqPc3BSz4GKMP2TIdo7nqTGNnS2vvkVepzfgL
IMcd8E41zEXdK6UFGRA6jXqajscNnKK56N/PpPQnGpbWF0JEz/DEZILz1/2pm3rNe42H5fYprEv0
5tWPeGsf3G/KAzPqlw/FObvyzgW6/b+cD2TBKgl3w2G/GU5WyEQNuPWMakmnrCeSFyLDMCrLD5GX
ubarFwEOGJAkdebVk3AthHj3ZJlIVznoNXNfQZmF4xjnEpsfTfP1vhd8UNh3ANWsS2L9wdemamID
UdhgmVNjCQ+0UA65fljDLXVqSgsLm42WrBJezmRR8e2mH9NosNyoSTHkYBYcZc/r16/fZcT7i0Fr
QuBK4w6vu/VqzF5pErLR+ok+8lCXhzYQcNq8x+/I9SZJ0fAMmVnYNKLiQMOwSZ87vm2RbdUFOvdu
jidEcNQUscH9l5QCN1aQSSjnu+TKGzlSa1nSYGdOLOGm8nUsqoI11zHJkX9UP1OEoLcco7afNyy2
BCdJhlR4HjxK54G1EAzJGVEV4UbIe8R7Hl5YHj76G4mniHiYvSW9PKNfcik5jsDDgLUTATyc7RIX
RU+9ggka4+Dejt6Bg36fgU8U9vb8xuPhmTBid2kY3vH1P2CPGQ6tnKN5bIxo/Wt4+/RDyxYyV156
ms6glaHRgyr27mTJwftS8BVjeNlFHUcSUtVP8qOMhsc42NypWA0XaV9zjTecoSKMP6GY722Obsml
F2FCA1FsjKak8Db3vte6191UqJ/ZEwDxzltiu+324gFryN6rJSkE+1eUIgE1T7r/IUjcuTXxX76G
wBDB8hFaG1hCWW6nubV8owQfDsFu3PJZu0egrzv0yPEfk+bqstaiYVmmSJkodPgNG5IBavuqFjvY
324B94XHpn0BrqvlJXXMzSktWRZU1/zSzPN1iGL49TGYhGrF/2qr5uG38RqjlilTvOVkC1B90yVr
sTwP4vBu8GVPxh66dVkde2okUjRUg9mt8vLuxEEeLsFmhuCkKCOkgEgg+9kzF05FBYRg+9uhfqMm
MK/4gjNgO4kCgRcGD8+nFrKCAN9UarIzuTEfKtB5isHnNA4D5b1xKqX7oSCbEM4H+RZSYtqKk1+m
IUIbcawbrmRc27xoZmkIpKbLARZE/1VWdu7nToCN3/0SnvJ3JQpNj92T2Br3sDwoYizFGrEvVVH0
QTjrWFt651GmHxgcj28NHwboG3ygXwIQ7avUV6Ato+WuU6PcVhuSB0syt5DJY2gSLxqwGLy103H3
ABBx2VApV3HWQucOtTELAH2Oo8chKpYIdTDvMimhWJsBve3HFclIyimbiy7m9ZqXP8nQFwT6OFI3
SUSBbVnFB8dZ8aDgDkoPx2UTEa4zh1tTSq5szrxDMAQlOmoXMnM0bbI6XmUvGC+cD7pTaXsn8YXv
+gfZUpLpYVjWeRJc41nUA/BiPmOjSHsOvTg8kKNlC4L8qYejjJbHKjWrqR+WRDQv/5wuxX9nTJEm
1fEvxS0PaRBwcpYFKbur3SEgjJw7ad9sAcpL3O9yNfe8qQUC9iLleMtwse5jQF6c5RcV9qVfUiA7
HrYu1yZ8sM1nZk6IlTq8O3+jclT/dPLGzRvfW/balkmphguKIMm1OaqJU+QCwTE0Ms+ungN+wYbq
mGHDGjm7OAPkq4cO93Wwj9y2u+anPfc9oQf0zTJkY/Pk5J8XzhdfkgpuGPYGG9C4ne7lCJQxcFlv
spUrAVURSR1j3PWAFeZa+M22eDHjhohrJZ0rEKNTeJEK1kMGn0WkynA1mcEJShVTznH91MvcU5/1
6u6Kv/3PYJj3rD0pCztEi4QZLwe9Evt55P14gqXMXZ26W2CpjqQTqvih0zp9O5gqrsS/+goFoEag
8G3aQVcOH9f8vuNvhu6prGRzVMlhAAHFUx4b+VUzP5INsI3c/VzoIC9tUusDZ8KevIQ4dBlKlNM6
zpABpLsS4/emVZaZMHvLR7e8UcVF/nzg+5GT6Z6x1/xT0ar64sQcAD1zRTxzJOPFU0bNv8OlCnj+
RQYwJ41gyrGhPwNq4sxukBWubPVdkbm6jKwgO3UAd3uuAMs+WrUwESot90RiETUftTUW6mvlN++n
MqLK7S0fGPfznpaCCwkKI0S5cgRNNNPRKFED5MudrPGlloON5digGaBJ891GO+dYOL5/WWcYJiB/
JBTJN82Hqp43Tul+/aanuJzUe1fGF0lZPclP6Wgf2p7p+Akk0cK+0krUeo1LaFZ/xXTuqTiMJD14
UDR9m/Qnv8rPRn+OAK/dXPHllkJyevxl4F58iyInFXXGQ5YzEetKibM+nd0d0p33J8N9ss2Dau+w
lw9XnnH01Oe+wdvD5dq63lv59XUhcRTX2Zf+GnTLs61cLUSWbvsBeezTicwz/i5ZRPYKV8tIeyN3
paQYl7aB5a0NIBVLvPBvcZ/iG+Cg6Gv3iSKiInJgtT7qNpa8cMvXs4a61ukpCf03eywe2jRKVUeu
6HOdP766duOaM3gaYpnH6TuZqRIXrPLI53aWNXabz7gMwGSQk2IRbaGQNkC7aZcaul0+RhBCtbG0
29QW/KGzS3197HjWF90xQ9Hoh5hXcUvDflxUEgS+8NKVeRIGUbiRodl6T6prmXSOqeQf7tIhig9t
+rZUxVaoDGhf6zB08thZFpomqqyrBBTK5EAiEpO68byyC2i1KRfLzvXoZoAAdi7ZR2Lmq/B4mHwf
ZvWj4TrECwNxezgiRVnb+ubvNTVoihht53f+34BVKlUYnv1xD+FccRNTtaA9/8MT4Pz8gPeQyDvF
qGxlhVZwnWdchQWm8DwdKsICrS+Fq7uujun6eTxYGJhRSut0db22hhcAJRYQW/TLdk7ZktlFaTGz
Bjs7TeBcigMHmHbL52JXabArhiRrUzuYwzzUP9CplAMOQ8R+ELXoHKHtcu5L9C55KkcmxR+9yCP4
qEjFLkqGJVaUcsUp1NTfcCNjoe/xmXyYvDBkync0Ube2eBU00VKK4EeCpMmGADk5DSiXRxkzU3Cf
9sRij3VTiZ4IK/+OqRgQdqYQj1XEUHTJUlxyXMfw2L+PICGOYgqgrCg53PS2rIJ/jwpAUCsTBQ9a
yg8qJaG9FBoXsvUyWJT/zcGIn9H4Wyga8IvM3VQ39J89LDBNcz661vMqMoLZMcqgXyHUh1cHoYz5
mdrM2xNTyTLiBS88SiIA+XKAhK5/5hIZA3RdBzDf0fRKKxQ4diEJmJlZE1+eWCLqNCg1LX4Dabq/
AvVtH78QOQEOg6wAYlYJdKNdAiXRba7welXqfngiaLDbIhXJJ0PBQ8CcNtJHsELjSmILu0/ix2bi
sfumXmc54P4eP1S0kyZ0XPplhLvMsobXDSSd6Ljlsepk42PHYoDT9IeHXZUybu3f44hHPKgTHfmU
JmikMpj3mdv+VaVJiAVXbqeM56XqJw3IFZPyc+xMem4chogJ0vGc/tacBCRXBOxRqYNvPLlHscP+
DZABNXwgcagcLxxwk8iC8ElUFrGdNjh3iuVFuEHvyC46z1sbCNx/Z0yyP+P2sfmsP7MKn9zDPdGX
Y54BZHlLbdmCprM1lS3O5Avrge5Fy05h+HqJ0BFNvL1CuZpLDQiOfRQO+nJOURUxLw9AkfCV55Ac
o5svrliOxKbX10alcFxAYKrZH8+rHlydII3iPZ6z2JMRyYolZU3qXwo4YFuEl8a/pYEtVr1ybsiU
NQyc9bCQs1gWli1WDXUaktpxCnrC3xOGoWW42VeEodT45lwRQ2tzQRbHficl8wE2vqPf8o/prXHL
s2dLp90jTgHUYe7ykI1diywHWtjySEsrmSjkbk2E/8Mj2pQZQSy4uwGqhWqR/tQdefwkf6nnfUXK
tXbwUXXUjq78p0MXUlI1APBSjeotHX0tzLykp0rfysoRBWh+msYsl219Q9vr5GeODY8ftsATUeJY
RRGkfJKQGBqtPJO77/fNxMbuMwgiiJMArSwCj66/tW7tufWJMjd+YSv9NjaciSHRGbSbuW7LL5nu
KRhUF5HD+oiEUnlelm8+EQ6Dq43if2EY/DIpPquqZhQBYBBRjzFDUHzkE+RJwFIYSZxT2aKWR+F3
ScF8pu5DUtXWJVUQaygiOqG8ysvJ64K8tviBQtnp6MbpbO0EPMjRxOO/hpW8qvwd23YTNAojz4kV
+G+Uivp7NCkFlxBefqEsAxzvcjZ7WyGShWFticv3VrdEQlFkDCFX2xi770fnyG+q/pJcRDSgQh7n
yaXXf7zl7DUaxhYDIVNimu+99IzQDNIxmGIjUeo7B6om4+z3wrykUDC1yzsT4GH6Sxqr6xH3pBFY
SzZvtwvs1rtso+1kl0aTQ4s57CuFwQJVVv+lZhDza4FpvwxDyPQgWZL7OD2J+Gwk2jgXQYQomATk
5DYebwkRGNjG9/35x2dPouzu3rpMY6c1iQMy4612w6y6iO92f09dkyBqtNI7KL+Zk+X3IGD/ebrt
kN5tjY5CCHTs128OGsGhd8Fe4j+2Q4i9+yc1i0oOzasHZMzwIyq6u3QKoWjrBgniyAJ5Qr45hgQP
cdhSZnLKxXY/bChZk0ASpeCpnTz3tO1JsaNlfh+YvijOC3DKyQn6flLiQzUP3GCgmHXbJWjebiSF
rSozUzGNoIRBMM2eKauTbWIp+wZLc3buQh5h92YPy+SfVL3MWPYgSt3GLzfJIU+Y8Hqx+LeqKcdy
Oxs07pWfGvovWo5yHFTgIbeQ4IA3PdhQ6LTPTuuZA3Pdfgym+gyiN0LnDIXtSm1X8ewA2wC/Urgx
7SvGFgDFVNPWRdf8+Zc1pv8zjOZEms/eKSX3Ybb/aw/JiP4uTJAsB/vvPJL0pKuUISwe/0M3ijoK
vl3s76r0/a3kVGCShLS5S26WhvQmPEQJotRC7m5mdsu7/DgzEdo9jsBmK2yZAwSjXfp5BkxBRU8q
YTw95GUKIp+5GeDcjlNrtF5xQ9iVAWXVDyAz947gWCLDKmdD61iKC7btBi1/dKpvEWa3EtAmHZio
OOSMqf66Rnkm7APA9IMfL3cG57OT6yemlwt3exKZk81bwyHGPjUOi+lXTltJSway9ZQl6skc0Uvj
XpBVAoPfO/lXDulit5aYW0+Oc9kmNnl8jBdWB8lPbUfX8Mn0c17qrZczsoMGYmRPq2hSiBIQ2y0+
s61RpxCJ4ACc+XXwvgl/Drkg+F5CSb2MqIYMUwdybyV9DW1Unuu4FuhcPpapLXlF5Muxo/46w6lT
s2t0KPur/D4IrbLQMZkVD3FNoyEyYQ9IkJaMyzUjYXZQ/gUXMr5FGme+U6y147SGkx03mcIqDAyc
y78w1DtrSLP8HBmbLYUsP1R7rV5W+w0q2aEedHmjbXW7OCJmJABo9TY0flYaLuLsvExS1KqwriAD
6vBAnhT02VClwyYQP9pofmXxtpKG/8Nm+uxXADUCmo40gfO2laTRtDMznj+Z6O/TuVVR1RMaEWOd
WvIYH05qcynJkCGcffZOedhjQxqAxNXiEk5+w41otqnJDgvhxcrkQ+o2Kla0FVNrKpWdVt3Nq+HG
QSQTkUM7U6VCaaDpcyOhc0sTBERHX/9MW96hjIFxNgWaEluxKz/28Drt7FcgMy/qhm16UD7plfO+
soGadtmwxIPj0PPd7z6URxYEyDVLZkUnAtQzuQR8JKWW+ZorCaunZoWqMIoczWrWRwWpJfpqF9uI
OEGRdn35iRSnSRtIhnEbvu0LKjNUPE9ybuRwYZakZjbOfqmhtpoEqcZ7YcP1ssixV0yAabVEnQOg
hWeBpF7RbCQGqZhcHGioZUOGq6Xp0aKAAEffHQT0CZ04mZCK7vwfBv5uiiw9XDLEcJMsiQ3HU9lX
/AxfKMMvigB8mDsTIway+U/NO/2i86eHetylOgZ6sbIe2J81W4OAkt8t3A2lo5HGNADyLwjVIzQb
mMhAm84ASa1dYMiHYepo+Wi86xoh91FVwpP0zG6QXPrdaffidlLwHuYhV7c2ObZ6LKO38K3NBLnZ
lG+xfIiVQBrfgnRiuAarKizOVs5wLJEzW30fhX77P2ptJOJM1G2A4RsqIUUSAruo95ctVZGMVHWo
cekVbmx35sNSbfJ7yO/WEtIKv4tUSvPcTqZa0xOVhObpTNFf8q6kuAEJw8Qq72puSeOpOZf5qw/8
1w81Tf0xf7YZntXoM+/Lf2n1t8jA4CVMYWZPuW0cDzXqvyn0Igf8M3jALjbdnFORTIWCdQoSGf+8
/bOsDJz3u5o64kTVCMZQd+X6yr4VEB0UvYSJTDCJlql0/wi5/3jzf0xWIyDVyVBBx8Ep9U2s7vK3
X+VtRtcXVdKxTCJBSNqPOGRCBoHAzJw8+xApsEG9yCezfRWQGv0Ds6lnBB5GAUP+tn+mB0t7FEH8
JljAXUohkS8xFskYf23ZjUVRjQu+OaqVL5g9hpLa9yXPzNn9Isx1YCY4Spv0CJqXOBAKXwco5tDl
bnZkZT9d1X1cGCOa2mU2otqgJfwtn7gMcgdmBpv+xe7+YoD4aB9dIAIvro3RqkgUHwofO1fjYQDp
CvLjQXPAl2PCRn4cwJJ5NH/3/EUlFpEOqaibpMT+zoOGLqN7yEl2VWTAGc7GGcl4JHylo/w9FFde
a8zi+yoh3ra6V1gh1MR5JsM8njM7W3cQ/GgibWoit8OzKfg0TpztZhCF78KlnqBiGhij61VvKbTe
zIPRIR/mVzTdn6MoPCPvEfIcnCF0iUeit9x4AsxRodWAUs73PMAQFXqe+dWl0HgPtWq5V+XSeh6R
g2YTtzQSiKze7AY3eSoWE5YH3djhLp7cOgXbGwXOlyySnaoo74d77hsvi9b3D2X2IISirH2KJeQX
qc40HUiWZULG5LWzq3W4qdfXutYyrFyl3Y3hhL/7c91ydDWp10U6LT1yJOzW4ILUaDRqH4f1VVTd
fiMdEn274vI1U/bSRTaI6NGXuOzf4jgWLAf2sM+rxKYfy8SKDzfEbI9u8cLKh3UHRsetR9e9pAHJ
a/i6XnRJVjbyoWPA9uQPGzy1FSwpvm5+U5+gZVv9LO5lJh76SX3KM8K48LWPld8pCcCq+ZNCdXvW
AmSCVt90OLSnr5zqo9MRp2vskvDO/P+MTxF6FMWouCy69qKLZCdfkCMUpaPnuNXOUwpUPbMqM0u9
G/vm11i2p9ps8WcTM1Wq1S+G3Oq8BuECLwMmaeetfEJT+2ZaW7qic5+sq8kJU6Fe32M2M937076J
vXqCVI3QLm33nXIWrKytaAaIZyLkNhKi6OQo2tj4xrM8i0CPfLbMsf1IbIMwMaF2ctcrg9ZGJWAe
cs+LNxNLCrgMNHpwR7mGHCqdKoIH7vQcdEGphs9LhVF/+S5DwUjWMaFgTK3erckPGmCTfDpjzzqt
eoHrXRs/9u0sco47p+Mhu/90lZ3uayP0nORNCSI03ENjxip9WCR1m/nslqBm/bj+uGmec7d5nAXI
tFCggXbcptsY97Iz4S94MaoCLrixklkSvfw0jO7yEIK5drvGDPMI6Z6mYuT9JWFFmu+/uAZ3nUnC
ANIwgk2i6uetsLgMl8pQgDn8BY6O6o/lDv/Zi2oeZFKB7p/asC5O+RoQkDgug4YqdE7mRmV3mwC9
1cyW5h0X2XJz/6HbqFqDkUnNUgZhnJbHKQdkKMxyh15JVGAJJxiCgywlO9NShhnDHS9mY1ZrvdxI
I1Z52rMe13HutdfJYY/3sI9fu0+D+L6Djj0gZAwK3uKE7UP+zYxT+sIjtOWrkFOj7405OSEIi6yv
XJOs7nfXxalgVNslMngkuvTIbpcgQB8jBaOzeZ/Q2CPI795CQxoKGCSL8IqErbAkPKKzINZWbyee
p+BGwVfh6FdUDWM5GvvIOZYRqeqd+XPH8ErFRPqn8Fz5OA3lM8Gfy6uRHPza9Y0Xx/95pqMFq9lG
AyA+ciWfAlBjqe7iV2HVu1cGAMWjQCnzKg2HW8216TyykI18UOVIUJhOviMJWwk8jtbAnk3HYr/3
C+sHcoPPK1UFmD64qtVOlFVbxfPNv5LU6ftfTnhvONV0gPdfaMOfoXOiY8I0tRbO0m5wZIoc+Iyf
HMAAOkRkSK1A5lvgiJwd2ZyYFDUyMNAxId1/GrjPWQgPExL8cASx0jaDiE9i08xCspuGi2IPsW5o
VUU2HQx1TkuBpuZOdQSPnLRck+pcr/tFbDjaUZmhq9V76ptSnLbUI0ld6YWVXMC5sGG7jOWD7Hqs
op+VtmAjRh/IEzZ1Pk1XBouF2erH3SSg++4w/R+mss7abgQW/7302zwLfc1yL2SsUFYbvx+DR5Sd
xCOGrtRFFei9xGBNC9Cpv+KcrZ2qmoLLt0q6UGjPhzJ4DYME4Sm95B4dogoBzC4uFb/4SMF1XWGJ
7zvL3Ci5xK0DFdQCx08rwiouUtNod2KEQCWgPqkSO6RmAdnsHWhZvq9cxNlu5OsJutG9sW5bDw8j
p6jtehddunFcd39af4JhWrRgFZydTJ3pfxf61XJFI1j2ntbpn0DE0CClZkfVvQ7ETyfwQ3H9wZlj
krnTotRU906vnYUTfULzJMdeTI2LWbDZu1DzAMzTOIQyYJDtGXwEkj4dnUSLvdH+EetZRGlkF6+p
kXdQSZqUER3msjIPDNAVrPxxXCmYLociLW+wABraSYlUCIndWQLFH2yVICnSW9BOm8N774aUxzqv
HVoR02z8FE/hxGla+t+ixMBiZFL1l6wWYl7I88JdYKhZyCJZ3emT0AEzehkn5I8Q870mPd4NGFqo
79lvtD31qm0rPIxgqImZ8u8IilVzCIlPfeXJqkgT6OBqswxXM4qQJge26cpiw4lhIYn+YPq1un1O
cV5lrMabW6uLfHeRamoXfn5FlGIz5wPkLWHlmF92IApFSvn1QPzhVvSggZGgYtiW2TGruR/0FbuB
BdwhlsNZsGE17mlEwcjJjxZMiBo+Yx0Oiv48gTosmSNjQ8O2mEVzQj+9Fc9T/Jwkb5Xtfk6/JIzr
365SAvM1hrzAxKraMdxIpDcusAStPdaxN0oX7YWJm6j+PmXI0IktFXuBmGEXUPV7Js4sXPsewbi1
1jQXPQ1K9rvNQu++Qh3SEn+lREVYHuWbj1VfNFOuszFQ7Admb59Dcmm69qwODkWaasRhKoHfRbiJ
yKI7YYVf7zGKnYC1SFeLzgcQNPhD+1MHsi+ooVtuhDLYVt/6qKw5XKqJWRIqX0QJM7dIEw5TLpaP
YSfHz738YKHft8vx7+DqEBZnO0efldktvvDqQMjfgjLUD0oWzZRsvFnULCXwoJK+KYeaaihW/OyM
8lXxrgJUG7C6E8mnLGpeFCIZIwgNuR9yz2LV0fgkLa175nGVZXKMiRz6TxV2vlKuLVLPsbf0vpbp
GyvgNvfTCBzoUeOSO9te7L55xe0mp6wrepNg9ajf/xP9Dq+91v9/zlhpmP+NW8XROuNpOEGpMwL7
NlFTYJzEP4t+9u3Ispn6cLMeJoAR53+ubJM0wnlnvXytZ+kZSBR+kbPB8d0bgK0483R2UdZi8jEl
UMwtKw7Nyc3cNDgaAYEAoJzhFIj3Voj9wJfKRmjOLmbeEAelZVLw3gxquZtX0O1aA2doPRFDEPQZ
nTSm0yfzeYboMMfZssa+f9uTEQ8JsGhmt0Ol6s/i9BYCA7XmpeCPEsvBdHBUyZdwjEOcuKv2YPbN
R1v4dSHrQo3L2Uty3cF94BiiNqE3QEsN8kd81LiXkdPSIQuMobyei6liXULZZcPe09TRuABSfQIp
REdGBW+aHeW0ToI8KGoyCHLh82LD7qpqbPnZO4bLyhxfUrimt0QTu6fTyHFieO01v1uDOgWaSt6p
feVE5kAN6JtwakffB9yTNiK2evWQR7LMixpmhtwHpNJlvX6HCTxiwu4MZZ5q14H+u09LcQMKCkb1
prlupGAKTqjJ3dj7grK/e6qRT70Vr19+h2TyWkqMCasNiWGqAy2/SsD9eMXimE+QG4p6IdH3d5WK
23vvd58y39bUbYpQsAQmwCqp339j+jWjmiV6IdjgXsY+X6EZXkFPB5nX6iGgoNTBK6net9uFX9eI
iFjmna//b6MtDBgA3Ya8/fnP6boZGj3QbN5i4m1xCBo4Rdy6wgpzsPweW2kzIpcwZuKEXbF2CqoU
3TTLJm89TBgQ7AYLgHWzNp11GLlanS8+ompk79AcAyh7xYFbR2KXp38L3nzMqXJcvLN2SAgcFxp4
c0hVn7+gLohHayTfLwlN4U7SobXsE6P/KHnKDIE9N+vaIGZo5Bex+VAIuZmHDp6waOBr0G1orsDN
SPEiFe7C9i1ejXTrHO/5tPuR/QHH1fudd+zRMzo/yr8yeXtjL2wO2AwfJFzjIrRy2NuvIoHjVddx
V4RsVn/h56+on2EkSS+HpNu2zApJAMDEGGI7Er68eu6M8yG1rfreW7wYd4sDKbASz0RmKB0kya0I
xq1kjex+t4MA0qJusd4e0PBj1n5BKCOrqJnI7MCXazbImOFjTC3A1bXw5DrpbQzonKjyATY2aR/x
IKnXZGk+Akv8rO52xkAskc/NPo8j3NlDVkc+SOkGR+l2vgrT4iNTbuda5XReJKSt9lac+m9nYq9l
VQXmjalPnwDOKxSixh4YT/ClS/uWJ6rIEbUlfbdrOmYwBDwyxbZjnLBauwriWCKq7910SGv/XKjW
Fml8APMmZdGvRVMGiKBUQjOyk3zMhj/ET5xYfTeTNWBekhL9ZOnLW76tWhKNpCkKpqT3xYLEj+Eu
RhYsfPhXq4xnwlg7bHEI8bCCixfwAHn9u9cMIipSjGioC2R+y2RjqWuxOGpdBDP9Qf81NrMPELwP
W+dlwexeJ381N2nQfdBvV/jlYWWNlGu95qQ4iteYonMPzJnEnQjV8naeRDueu45OKiv8YVLPxIvy
i5ZB3voQj4/xugHfbG9MKCIjsZaIZps0fcwoS41uq+16UWLaMKSiS+BMfFeqA4M3zen4OIk3UQ8U
FwaQHxsvSCqUgvVChJyvBQbDHVf6RPtwqBFC+yAg9lacOps5EDj8TkwXKQ/rWee0gnVjFZHmhj6Y
hzM0Rj4HkTK2prwOKxGdMFin6xks6EMF9E/SEne99XCrIu4eMUQpQwjSWyOcVfnpUrJrEMagAmkB
H1qrIK1wsN1Dw5ZzfgZkpwKAYHR3On003d6ZHl8jjE65eidslDNFSmm5Zj+NoDjY8I4qThGOAqSj
zCJUFldXZ6JNgW76jJsuAyLbgpKOsS1z3ts+9cYDG2z2FWQol3JS2vTzkQVU7DdcQLR1qvO4Rp17
id63HMOI5xVP1RJUdd1iixO/nmaErOcaBa8dAA8BRpoS/qV4eW2LElbHDQ9Or1P3cgCETtwhySaq
FWiG8MuvZ4qBX3emo3cXYdK2O9HwSRCqHmCTexCzi3bcKCR8/w+NfyC8x4OuzU74xdBM6NKpDV8c
W2Nikvf6v8aqDNCCZpT5qfS0qL4eRq+bC+nQpouqWu844GmuGFi/J92Wfj7m8eVCJs53C6TNbehd
fWbgdhZnrm87lWhIVcLntLxUOil/FjB/oYt4vc+oK0FCcIcWrdxFWtk177h75BVGBN09eQ2bTXlj
LoDgyAvw0tZUb1/s0/S2AwSNXOZu6L+cKJx4ZYQck7zxZaSwRKMfKgwoPiJ17absvIZPANWBZK6G
Gu0WmphdMTUtJwNrJauheYs3heQ/gie4RfRKVz926qtBCU/uRBCHWp/cpetuH0mtPF1CRY9O9BPi
V4x4DW1lGeGIIj/tlTJRPl8IfKxOY2MKF1Ypr1yeyvvWGhMnw7mt/0bxEelYPQCjZtsSYfCx7lEC
ybtNtjq2Tc6vdsghcvJIcewhCgG9b8oVDtS9QX6vi7Sgs5fyVq7ehFQIv8m1vqH8SZSGZaZHLBgd
to4/7uH1R1T3ToKJeY/LN8WDqfF4N1KRsIIpFAV0RYbTzvWc79FQDfWEU2jdkctezsgTU0GHBV5t
d/zbMxendbIeGs9MFZZ2A+nwua1A6rZeV3siu2toNxfsEiB+HOvDQ13B/PkXre22geNLv/HBATe0
HtpTFHtJTXEua29JjCF0Ieg85Az/roAMT1t9fKfw2OWfqnH7dKigNGOfjd8NTCRkpFreh/oMebrm
foBC6/jjulMCfqsyXvLpignhv0gDcxc/TLNbku82FM8kl8VOObqbTvsbQ7rr56nRLTP/bLlWxPbm
ngmwyhh1Zo3Fu5IefacTycvehepfbUI3jUARl8jFNC7G4aKJH42cAeFVrdxHJ01kqeL5Pwsopnc3
msQNzZgGb8WEEabfAdnqz5XXoImV+QR3tNyQgeQR0bC6S/ehtvIcVVHLFuwJK/ubHRMprJ8fMWZT
Cnar46TjzEk8vPcJZLYVy8ewY/TazVmzV09BLsW4nuvO55/JyB+TqV4Uydt/ashr1Np/sN+i+3nK
xzv02R+a2395SauJoNpg9SZ3S6vvhQVQY9UcLyTSkGL4zsiN9GyDUFy9hy1SZNzzHHnkqmWIZ2JP
2tT9HijLJ1/u/nlP/sCqx6gQb/mk2JsRXJQWJm0gsllZX0X3ugCLkgJr3yYxrVzd+YU7jShzpa8W
zhOSponeslS8jzmXDxugh7foVPjuOPpORQ4j9soB5+lHuKEGk+clcJfNJnD3jgoQNn5hjN/NqD/o
WzmUtunqqwCyl5wxv3EOvZ0Opczfa0+Hllm/UrjTeMsRpunkh9ks6iGy7f2RqXdHTkF4mlDd3LY9
0ykgXejJ5XG4AGOMKghajIyzfdj+I4OE4wuvRfTYdg1hyRz51dmN7yszFL3M6i8FjvX35qIgeCh9
8yB9eJ0kQ5E4Fy7Dw7tGTKd7g9IkkM/N3I7M1RVtC9BX7njAuIYGypbFFpcpVJJemmRGzwoU5n9y
+P645zxuR8ywK6u07a+LUG6p4KQQlmuPsG24Yp/CZQ/UzcY1Hrbne54THiRcfYZFKWEYcT3dAWOx
cdshxpRpv4WiBkrkRVvghJsFu7wBBJfrbH2Z0h4nLVhzF2y3IhxcvmpehtrZqxFwJYFtnsa2Ib3C
RBABnOEgC6nCPk5sWys9p8G/pgm1NLXY1XglWzPkxrCJQ+/q4JMqyURt7ehFB7f1c7+80jG3/p0F
Uec3IZ0TN4rTdklCP8VwTwc3C/4fXM4D6DmjoDZ0coTblY2c0dzhJfrcetryL9cKvFEBuZxKBeFe
fJC65ZZ636iynanrF2o17k3OSda36IV3vmygxkoNGi816bQ1ZeonxfVcspVa+1MAhRTYEFiC/mKl
tcSzRSXEQZhr2RDJWX/h28BjKK9svPh8Zghc91sGuRe4uXOSOflHsApwkPw3RKaMr1SJa/qQ/nD+
542W6liNsxWtWalXl12WBLY9w+YkR1Ft24mk4Ss+i0XjDB5lZqdDSk3XZFA58bmYoZ73T7ss0L1L
BzpoTsL3gcGGGzc6Z3SfSEKNP5UzbdevXZRpV7Sn/JIfMdu8F3Q8Pkl55q8vvYbqzV5xDVefFufj
IN1dD8n3ulcW929oGkv4CGDLjQb84vAGecpjNLcCUdaEa2knK9xNDglcGburmS49Tj4+OFdakz5w
e5n+32DFITOV/Lv7tyl1QWCpwchnOAMr8eyvAJuJSI14O2wJwC4ET6adb85DtCPh6fZ3xeeIQI5e
59Z2tWzLT7rxy71/IE784Ha+5dtCT4gfBxn35+qOTnJdDeBJ/WQ6fpZCfwHMsosVcasDizV+/kyn
8NtFWbKjq+6E7tJsevQamkLrIQMYzHzIYDEUYPWL/Hs+AGnEY2PodbIyWMqXC+GPmQnbxdJEe9EZ
vRwiKK41JhS443WuicXP4rJm9MKy+1WG6SFI8RuflbetImBcpKAxOnPS0gUmcI0FF+Fra1Cq/g5Z
oTdWiY2o+fMze3fQtSbwIWMhGcJ46qkvb3qyyyJA1OPR/0xySvZ2/b/X5bDY5TbzwlEeoU7sHFPB
fx1fP0Tw5GaNW0cjeSJ6Kz5qZHsbtTrUvje83JLtB5E6oXco2UrxidwPd1r1bkalDUwtE46V2RAd
20hRLYXMfoF+ff+xhIuw2mp7/dSTgl9Sj++9ik8J0tEsxD3yL8XZm+LUpnnL9tUmOQL6O1JqVjsG
FQmq08S82dXjBK1Us0elsLgKvzaKgOxntv9f8Lf5M0TRgngSDRwphbyUqkKL+k8SYhSqUAvFL/G5
HLzam9VxvChLon33ec5xOnlxWcdDDjtBadjIG/y9W7XmWyRiPPGuwA/MxNnyy6V++yShjNV7Q7xV
3QSBIc1JRPpCo9JByyT2Vzwcptm20tGRAPX3DTTzn6DDCEEZeGp3hB+qRn0ToWpcjSsSvZxW/o4r
Du0VLjrEZZhmaZ01+4ClBCeQJASCNzg3FCA2lkNyOwY+J7Sg2UhELsi/nFTmQ6kRbDHMaBDX8iwh
OcPFxXvLxlHjERJGvYNmq4txdF9Ts3mOwfPzZzhmW1/s+f90w5R7oWllbuzTJaUq10BgpOS9bDTj
koQxIXSHhAhVNtLk1x3EE/uvDHHFJIFU6FnPFYrtnh46U0ZIUJJineUxyHnMhBplA+T1VHR29MbM
DWN3uqJpiIGnfs0Elu/g9d9SvSBmWs75pRJ3C2z4DwxAQw6X5S2B67wiU2gJ8InCRlR6j4OaPj/Z
cDd4G1Zb75F7c0FEWyCUgE8nX1dFDrUMjVdVt7SqVGfL7/e1d8OikA5nfjJbfA4FYPL6A+O3rR6b
yC7dRJpL7ZW0gI1cusShspb3QnL07zp+m9xKC8EHMI5/zoi6ieaSw3+jqbEnGFQZr4x9sC11XX2A
udMryxIp79VHvf55PLlKCsRlpTYQtPcsNqGqHuELsG3bI03xaeYdsGPvr7lyQmNpnIp+WJqvMhxu
oyWszAvREsYnueloWD3PPj++Zat3gFjU2hpXNswJN7mK5J0pVG8UEDYEqUSZVJOTchvz1qnR4oGX
gBvHG/G36vKS44aYSXTibhq01TQ9i3W3mqMI1UXnQy8ILjSEpq1kNyDw8qXtzd7ZS2vGA8zxd2un
DLbV3Glt6SDDdemJalWBmJp7pw0ozuJXYYiGcCP3ib7/ycJ3gD3OsE+jxSS5/sgvlj7fmwR5SH+m
BtH/qnkIAmyTzOGjPKTCgPy4KoFwF3iPBe1XjozFYaCQcKsos5EmYfmrXVeXfusgxCITvYG4CRSc
VCF6YsLaTE1/yd5SiWC1xOn6WQqTzzDCC59ACdwAKUallgnSx5C8abTxFdm+UalAhmgDm9in3Utn
IlLYq0MGxUJHeWWc3cz9ANnOfPlbhf2iN52r7hMsbmY0Hz4y5kZNwMypEOo7k1PGq4Tb/5ltIOLl
YCiBtzAevgTNJjnhApEKkLUYYa8FNlea5tNxFTqJ4blX6QZZT7yYwUundk/ysK5U2DjvPs5BdbWH
iHr1DvwRAWMpYMuqigzq8C6MHY3hC4yGHyZFaZCrBj0fPT92E2RI+vWXImFJGkfF4Gz/MT1gKwK8
iUltia6VXVMEvLPWNrRf1FrrX+J0tMJ7hloUpneBkBKG90Fllg2a/gXiGYJq7aoaqElt1tGvmf+E
Q2+g2HUoOWu9/ugrY3fGbutHRPUKvlsawVrLppdptqxZjdYqkQ1oTcBvJANqrj/MBbmVFe3L2nfc
+E+mGDFcXx0IsxnIYVd5hNWiSmk+EOg+bVORI38lH2QkSAo/gqZS+1oXJzaYKxY8U6WzQ3bqo6e+
32aNr3wAxIM+dmFv2FR9OuSXDjPDwa4CAmqcfD6izNFDlTjARJHAds5BnMsdlhuqInVGGfCubIwR
7cB6JuHHdZ0UorbVj9zn+iqju1kMVT6AcGIhXXtrwaq1G5YyQEHYvhKpX0mhVjtIAyawpkR03ZI+
TlIvqru3gxmD3xK/9+cgGD3gAk6vkVKqTZvlKQme+LLAmrjU8nWd/am0f6kUrCWXqfIhfA/FaIKp
VVcAYqqimrdRsGM+8/5EtdV7MAn/Kci3CUZ5a9DE7qOin+8tav/2XvepYFrj9/lwJohK5E0OYDzR
FrAQnkQrj9Ms5Dn0Gy2JBkq9yswG2Zc9gbQg5D9nIfDNlncKD2RMuu4TnA7sttozxxNC9wt9Jlvs
Ze67YD6rbkB/Uwxlew+0GQ/3PyWLvhdz4VKSKICq2mHe0w1EDYP6vpKLzZGmHHX9cCZ+zyf8tZ02
tJ81nC/ppRfGuspxb40eBl6+hwDGZ9sy8ZwXilqOQomgHyaVk1Vdbi/5IelRNWba1n6DVPPqPnq3
5/x+TWPVbGi5vxjPqVRk0eWuiH+UaQpBxbEr7xTu+rbhATN914OwLcYsVF9BIiVdFUC80q8u2jah
uVQmL23yVH7lDRidnE0D8w25yclYXNTA16uA82GKIGw17I1O198ZLroPwncwCpnVyjfNANFNHfqp
W9g/tE5ULUT/GUc3z85KtNx8BZdF4AtNbEHNr/ayH76QriDiUCfrkuRaZjH6bOS7Gs0YWGxBeTYa
U6+QuXllelxRI5tEypwAM8GAg8Lk802Dp4ITemrnMtq32BqUJC9uBiz/PjhwPAVXcQ5aBS/Q7GNq
XH1N6fXnHEffBmHsv7npLEGc6NGYZTEcvoYcZcyr1n+yirl4lUYR5nFgKo+wDTE493exRjOX6NYS
I5pCdPqSO4WnYg2T6/VeyjVCjEibLfnphzb3JYOWmg3ZLOe0uP5F27tqsTLZknELHvKNXGJfXD/K
M5eHVSZb8rJrjmNjK5qGK9XhEC/CCSAEtmXPw7OmV3l0dT9tGSbUF9zNn25qMDIgf+Vym083qz8j
NpBOPjjTWsLF0PogjKphchmf9TO5WOfIhJRMSdOJLvyxUJMyhU5O1kYWsOY2qh9YaYPaIJesiGEB
8oMrFPIiM8+b+BRWJPvhBOc9GWXwf16ydWFN3utc2X+VCUa1CoqIwBFj1CBeTAUFOY0JTgDHR/IX
Ssbv888eXncvxth+ng/kyt9AAdzGUQZiGDMrX1t4Wtk9OPADGfsw2utLRzeu+us8tLl4hotNXsQg
XZtHVVYKZd+qh7YlrLj6eEyHEuwvgSt6XMFVzbhfe7/JBJ+es74DqnwOuyVHMhG5jcgwrn3bBpaX
j26EkosCXg0FKxxWK1RqRpT7bCdo3QWdu7g0JDRsqTK0ZazKu2p4FCVH7jVsYJRNWmRr3Is/ZTJC
kjVU7gM3ffpAvjT+Vb/l3lEmURrOC+niUtOyNiiuuzta5S+JqAnDKS7RRTnHYonFf0/Z6gmqEfTW
WOkkztEq76wYBL+6Rz1aclu4zRbEL4XL23pJ+npto2LfIgXsu5qQOLbrvKE5wo0SUnqOh2l51W1J
8zdMUkNJ4JUzKo6t02YvRgsU/zVK3Dxft8/39nBFPXpLilR4pmYXZEfV3PUB/Ys0wIQ9E6ezWbN4
0UPuanOOU3He+vyeG5wmfQvOTGQO8DQNeU8UAhv+7f417x43MiCs/yUQuss93tPl5O52O9+AJEgz
LANtcuqwD1Uz6nww3VpiYRI7h0uynO135ZjXog9lT5mbnxHiqjA+LoXF2yENWaTPAumVXDLyMeo2
IpJKAq4jF7jzGMGeMEbv73SA2wQ/iMMcjtzwPncJmwp0V/WMgxVLPI0HIEZh8kgr4s1yOqVzBwqU
Q5eau8XENWImptqmNsv3JxXezMedW3mCuJU2Ox2T5Twxu5GCeO/tPnIfcSxP3KHk31uamcqFXfZE
ZTQysikqNlQ+sCOXsWyMbNBUiSFh+GfCYQoGwO+DYW/eKFZUzjHeF9olbWU/puedTseSbjhG6jSb
N8pEGTwzp1KPH2aD4hDCkp/eDuvplk63OXqgxTcbHHqgfZ5L4Pcc9+3uNxCNLNOpT7/WtxeQgnAx
kZFEnFhzkzt0FjI5Xw+YcVH61fP3elAfY0VaaGdqPm6iYiNoyCnL4xrB9Jjqaeaa3GDfrCbNvu9H
XE5WCGhS+UPQzhZBgbHUzjYktRjZEEv5/YZWBLB9SFIc4pi6JoiCzUvifyOQz1Qifvh97Z1wLBXH
5VkS79PIn1MA9w2c1o3fRt/3C3hShHIomojdNdCcFEL8ctdN8z8/Pd4lXs4cNGqJM84ybIrV2at/
KS8HdKAKblk4b2URmaPZMPmUUAdRu/eEdUaXm2BG5SrmWENuR5i5jIeQlHOijhm7GuMHN4WFv6q3
SvcSqloJ68ToOJkUF1UD96t8WwJBSR2C98Yyh10VgSGtc81FZJrbCMFJd1iv5JbASd9dnm41khpn
i3Jdq7/7Yzxhj28OfsIlQeWFnPV0w7luI/BCcg3Tc3pKQWNP4YIH1LDXrJOLis4K8Hp1hNGspBTA
j4hBdyZBOy/5KgUnj3RN8U0mRzmPfTVqb/9NGzWpmCrb3oOER+jEwt3AOnJi6mcrrLynGaQRCO26
vNKJX9UoCyTT8NVlaHZUYHsVKgtn3Az+ptyO+ooaW7nM2Z1wA3UJunosjv3coixgwjQ2gxWK+afT
d4hwkpZJWCKUKdBvpHnHQaRrfmScdIikrVuH0tOM4I3F9dAZ9rUc1GTPTy8VqU0yyB5i0oEZkraL
AHnrWCNBeRF6LTT82wHEV9/8+uU54MbkHhBUrpu0TvENFE3k7WW0UXzcF9nLJQ2y+XGCbWlfW7iZ
dErog8VXUaHncvyVuog4RKr6g6bLfL5Fp+fqxcUAmUPmrhvf0pnfj23/llN7b7ozWbEOgr8uc4jU
UdY0TUGtj+yUFizVNJrMfGk6TOvAk2AVK8uwuCyBNePZhe/HvK5JA4Dqspkv5gbqfoJQYxWUOWPv
0cZ5tH2RgNJuZRCPyQFdqew2JZ8O+LSNMWQnQ4BTUGBy3aWEf+MeICUM7RM8BCLefJaYqZr57FG1
5AMc+TM1FNeTXxqCvuFVhExgMjFQtKZoRnEG9uZQxt+8TkDgSxN8b87CxoonW4mgFQ0EcWiIENmd
Zsa19WF7yBkvD1eM2ftZiuH+CJ0Fu+ljagYzVS2NZWzzNlwDI8dlutWT1e6E5R4RAuegIWsiLMN+
arDCEOzePNuc0S35lqyoIB6v2W/zC2BYVPeRSF0y5mp/zqNLBrjD1BIYpP1LhP2xCzNqwwrA+9/t
8MiLM/8iZhNsHu641kZ4sp6LNTJbt4q6J5hSx/z2ODC0tHOY4CIjRJuVZUobArDyLEwBEzdzljtO
mjAlUOYE/xo/HXcm23jMcSAPURjZHc2+b5QnX6fuEAduWlwVnHO7aGlUFGK4gAJqqTVr0oGQ29ma
RiyFbdr1EkyxQQCRo7NKBB6K2IvwqkzRNUdg7IAfmAuKolUYoGSJU/YAXujCNtkLhv0Xp7w5xMOV
YQ1eUSANvpZtxIULU5Gqnte5O6CwQG0beqGmu9lnqOi6Y2GR4Y2hhf6OAY27lPDknCJz8R6NIAQV
HY7Gc2EG/xYBtfwu5Di2wJNjxP5EM4VM2+ulGgw06ijwl3F+tOjf+XpSgqK9m4tH3vUr8xKYHnfo
hZZ7oa5n8A+AarEKFo5qnSG69esWr+enxCAkFMxmn6VKfUQQztIHvicryc1DatKp6B9EUVy3VIxd
4olw2UZcK/Tx6+qtJ/5j1G/K6/EqGdxJ65ujduveMYZiMThSYHBtBKZ37DspDCk2xu0Ut0GLMxiU
mnqAiX+ll3xBoNQigwOF0IOSgBGbVh1vGEFzMJ7EwPAA8zCaEXqqVi/pLBTROo5gYl3ryGKjuSrJ
pSMlNaiY4Vt/3srqeCOdLBKJak69VNzPM0007LtwT3DwIYfmLxLOhyrOKfr/98RaUAoHO2UBa5xf
9r2s4APYZkAtkRXVSNz4eI8saziakxPx4jVdFuw82OJsnjPdeqmz+dND5zeAusHLLfvAH2K7TrfL
wnJLTDz7zw3fAi0p8EZBBp7rAjfvxv4xh2FJFiyxAvXtiMcM4W0ms7/CAvl97BMB3Anm+JfrQXRG
paUxHCc2KqiugVxXD24REy+4j6W9ybHYFOjWLBDzcviZgAJhQ/F1tYEX7sP2CTN2Mpw5Q/B8H0mz
6KsgwVBnm6NeBW8J3oSFCXOuZ3L2vfrFMHbHt9nTfEbvMflk4luSupm6y95pp9Z7PBsuCnGf3Ph1
Zt4B/ta+O4WHO2otwCEO87c32/91Wgll63SSmt/Aoa64C/8oq0hwmjsRiNoxqbVNX2YdTG2+2Czg
2zq7JSA8B50G3B2CpGRHWWSTiUdeMkXwFLVwsT73EHp8+0ovxIYOAfTH3dyF5MMmf4LJzF6FKiyc
0+Q0mgk2oh51r5tSIG6nEdu4j2f3v+CG/LBYFjmLQYYvUIj1CJ+pfPWCGYTHLwUhml6qf5Ia3ZV5
nAveWh+dk6N+Q2U+V8yRmRbTBY1Dn/DbJc8taVr6z2I7dh6SZV7gThApKX9B1qQK32YlvbfbtyN3
OOL92I3GAZg1GJmWoN9WG2nmz+k/HhE9JKT66e3sRX0KOA10fUKAVYeYQxpR2iQyaLBOtQgM9UlX
YniJMaRWXqdi3jbgQfyCfrzm4qliR4S8NJCCf8GTL+NZDBPzlne3Ac2S9M9sx+SOYlmDGiME5l/Q
4Y2b7Qdpd2gDQ73GHm7NRAjKLnh8jAeoY57SiBbOhzmS3HPyeP99eeq1z2aqDInz3rAFVNjdkl/i
2Omx5OybgtnL/nVBXW92WZ+gTdnng/n8gHgpD9XjG0cU0aOn2ILsxd8Sr2YBx/DFqeFDaMVyY4q6
Kz+Nlv3g8ns8eu0mqBEgv+98dWch42VKlFFoprdxP3Q2rDcqQPTXKyka5vt8OK0WgeLalXaJS/35
FkYjmTqPisrbTujlsX2AtYW0YcAbY0PfqS/LWtFAI2E1pQ8dkX7jP6dQUFfblwhhG8JY/Ehh9YHX
LsH+0b7Fax4PlTynJ1mbyrzv+Bbx622NnsxYLFEQ1Te9tFNHTQpAiZfutPB8J9WUtEBnyVpRdjmT
LAHC8C71QmjWrGyLB050Q/kAJRXNNuMgVb004VgdM9RkeeQH07/KvzRx/n4/SM0qIdM0ETQlwwJi
fUYhFD+cJLbZ79/3oTL0VE7hilZ22890pOU+ynMH15zeivewLrFkNoCoVax3Ruq5/q03k93mZjBE
H0uOcJl29Z8cCb9yIr0t74ihf0KpC74YAz30sy7VkTjFc2IA8r0KuF4V9BGqYpr6gP/N41mfPSbW
JrrZALNjrI9eB1GT4ztmhEkP8ToNQiQ1G+lEYU6yMV7T9jm4ClTMgXG0xRG0ExQCWPr3RtlU1Qxf
wzHXfy9Vkn9LBAqlVQvDzzwosrXEUS4MsJlNCpt2DgsnvqjAUcx4eVyCfAoG3whDN50PbWk04T5a
k6txpCm+c3ofMb346zcfQyUBnV1trOqNMezJ+DoXi7udK6WKwZus8f8ceItW8LWoGjd5IG4eYTyD
I51wlEvGGZyh6jR8wU1YSVy/FCb0wi+rZgD8s30LB5KBkdyg6rSbhltzLO/PwvedNy1XLmSaeM5G
jySRQP4Glowd511162xuhljwhlePGdC5zbSHTk1+/xg4z0OjvtvYQqFSobVpHu9mqYOPl3bb7LDu
+nAK4+rNSbqD45+QASuxpjY2aHNWI8A653jhWRGZ5N1MQCvQxvODn+X71Zi3hkiNNN+ohFt5dJJe
kFt8Erz7SCWWSHms/rhAMesjRB/Mnm8FLxT6bwD6n9hnUs8GsUQ2T7Iql1fLaU+OT3J4zGKFGfIP
urlOi+TQ0D6/RQAFBWmz74qDy+WQ+u97ohfS1Z7A61X2CIu5fBAKQ+CQbPaxjVz+ijBIK2qZhDvJ
EnKSkfiueMaoEfpcuFs6zXqhlksNonW8XURkz0cVKXSInia/e8avm5RWFhHumziHZbpcIjaubl/m
dAfHkeIMHGbBazNkq03cYyroTGQ2rUt8D8R9a7pHC732KVZqObwUQG3Dg4DpPZ0kz24oOFMM/6d6
qFcYDc4rBGw28dvWRULaptslRQLJg1IL1RYAEGcObgsQIf1GJYyBIGzT1ljdmtelOzRxaE9B6+SG
pUUglJI5oQarvICEUtDci6JXvKGosUcTgtblhjA8GzpylLR5NPFmjvkQvVxYuto4GqpUbtpqE/at
ete+f4nXRfHD/9nq8HEy0y3PWi5v7PRbSr+7mH29DBvaqgaA3PDmwFPgn1xyinMTKIlRd55q1ekK
m4afgINF4LBewJiNkns7lp09TnDbWBM78rT9MUUheP0sPfNR8JpQbGKoOGHsjbQGJ0PG7kzauDez
YcE5tjOGfFZDUDDjIZljErIu7jpQJhwU8Qn9T+oWp8A0u95bSzm7LJBe47cARqhs7quuTYMu/R3z
Rtuwq5AI8yPiwiAcf7XxTI5XkgmQVbNKeY7QlgYVpnP1UAUEGMMUl+/LHqBa8wO8QspZtKEoKzG0
IFUUxRpQ0UTQakwnYziso1shY1lbnmf5A29Hwqm82mGRL6UtGqUXVSdi75vFM9vG0d6vM7kYEeNV
kKJqrvZzf+aiZ+jCVcn+FcB48VEClQSC2lWo4fD9T8FhRh7EuM7pmWRqbXCzE6hDgqZRK2Z9fnnD
0lkZGCCMKkXBlfHN9v8b2Cj7F60EwTh9MYdhvHGZZuxSB4v+2Jc8PYee+96MPy2lXS1SODTD/1Co
hi369bJDxBJNwzTGX3OfJMuG9OU3pZe8y4dZ0D7X/a5QfIpwZqmoRo43BHt6PWeFmvk9sBlR2i9Q
7gJGrBgKlyI47HAW/26sc6/LvDGYnhQNIdUps2SPPH1Sh84birs05DP6pJ5vrPOYGjL5Rf+Z5/FG
94ih+8pmvmUxwzP96q5n/KmYVymbdL5VsI+yk1L1Vyy6p2uT2HmqWSFm61OLhLsAgknMY4MLdsd0
b20KzREzHOrZivqb9ZIGx4L3yeh0yo0mfCMcTOatRTSDn9iPZxtMyzCRSXjQNT5M7KZwjqczza3M
l1sqUrqdWjF1jXFaoWG0XdNYeccA0Oz+Sv1/G9weYFpWFvJ3pZAKBj7mGYodfdWpshHdXjVjPPWn
5j5PcU/eXGUy/1VU+TV+Uv6eJrwF7hNkC5uCnOe5HiUn8OXOUGgIm3bN0NTVEfNZ7T5ufpvRfjI9
BA3GfNH0LlPSGBVE93Qz++Ei0vr/ORWlS5x6zrbpU8xf1Swx3btCRxMyUPmagVKs3f+5Sooj+cSd
kyhfwuil9KF8t+QGqDevIAa5zEf0C3r9scbCza8TRDG/dakwi2khnOipdqOh+femVPqqjfB6owuD
5D3h3FlCjS6ZK+ctpsYc/J1gjiXpgy9+ItrY/GAuIs/TzLmlz4xAdoPR0qa7cUcGZiz4yo4Pe5yt
x3Hfoe3sqEEBAtT9hqjpncAOgnmEQHRcbtuZTSJ2md1SYf4WWzBCgfCETHTiIPxzPhGKmhG3RGZg
Fhp0zslVTMRK51k2fdcWHNfpY85HMJMcCZEKn4ziY9MdRzhA+Pn0UqYsGos3bOmTCtTOb7vTWbCe
QeN3G2UrZ0B6StYtXi/rbymD2z9yslAXqTWDBdCVK6dNaV8zZn/hBNluVohcDJI+194v7iRcjaxp
HyoDfOrJ4Y05vWDTOAApnpO7BeX/OfLqvXgaGviyyGR4wqoQHTyErzZH+V2Nrnk3EySKmiUFflZx
a3h7FDVDsW44NiyKIrVoMs2xZ2JuXPgw5i0GiLLgppksTty6XQdq/Z33yxX6UCxEgtK1xQl5xGbI
GFqJixQnnT86JFPfomiZAMNMW+3Ss5Q9mb9O1h7FazFEoBqFRo1zDGj7pChxOehVjqM2+1oN3ad7
m1CVK3HXX93TKuQbT0Ky4LQfdJS72iJqfD9HSeG3LQR3erLeHQa5JCkZE1X2KlsMGbC5B6NR3Te4
GmYTT//nBaTplyGIQb2XSN+eOwmgoK/e6+dt1Xj8INSNq9xktPR0xnArZNVXI05cQtLpMVrzXOpD
D+7+CaAkK+GVqtzAeUCCB8uMuVvq4V+ypef0V3F1cvXXtPcKUDLpNIFxHz/WxUJ/3s2T0O/EL01O
7FACnObIDtX7TbmB3NtUmwc/tRP17ZG+FwuQFYnbIOlFabH1DWcj1PLTs6dIiMjgNLOWICTNLzBi
syHyfd8el+RXpvCIDHJR3j68MWqEoTK+TEk4kXvkL2qUaE38QSizIeI8rByV4G8kbOTsWCARIp/S
lcDLW+/ln5UEbDgZKAzhu9KkvHe2ATDQcEIV2ZK4MAaBBefLOjLpoPfVNxvOD2RDdjqKBbwF/2rw
b5eEGMde1BpcgAZdiLjzbIxO5D5y8Y6GQJMkyud1eTAxu1+oV+yGUnCwaoPVM/igryOntH0ByXB8
WCwalRL7XM1WGZMBZEUChqJyjUOXksfxdVrfE+r5DUa6k95Ucyp3ckOlKnUqlBlttKl4WvqcOBjO
Z1mVQ3dXjFdJEg65Nx2FL8ej+e7QtX4BCP2Zpu2SrOFlL5VHWQ02myHBmdmqoqHSznqpwT6RjA7p
af0CjJvafD6XdztIADp5WINAWZnqEYELLxl1HjfG4GVzVaqybxawRENCDGUYglEDO4BQ+8g4Dtgk
UjkWVDeb7dvhKeim/NYAODDN7n/6FsWfsKJM4hM/kIcLOQB+rZUSMl6/Wfy2oy19HtT9qjXnFnTq
pAXHwjtoSTx0M3zBcv6CpVlxKsZiuv8ToAxgAZmKLtOeArGzUDFs61gxczcqjHCYx/29Cft7Euw6
E2zGUpqo4tGmrsahfaEd2wSllZ/POiKsVt54gtpz2EzZCM7tqGuo9/VkFoievY+6wy72axZYPP8x
n5HtWhnZbUC6F9eGn4oO7xBMvUzNaHEbvEgKhJMEWNWHMa8dAkCpj/aIQPqi6vYPndjV6pUMpJC3
rwjZkiT/qP8NFd2HXT3bBsVB++nowD2ECBUMBlnkyaitGXXmncEKcFfHc6bH6sSNxKl2VSYqg2m9
TvxI64O7yG+XGjNWTGRs7tAmtDw7eqjb17EHireQbfI+qyxLCRoaAtS8HS74ZNmVzsSG326I1zKi
0NpyoeI83GJryRa12bhNN836GAivKENElyuIXgcIl3mwhz05/buevle+2r80AR2S7QJAdQXmwIA4
GloEMKMC18i95RizQtD0O0mjhQEbsVWHujo+XCK6Irj3rvJr2XSLfSbWR/t0B3dSQ5L17i/tCkNH
Y82SwMExCqYvT01SodXrxJnnNM0lgUJSZR/Ux9Hglf5HR2tukNaQm0W89wAkXq266Romxi5fzscb
tRRNzyRp/CmNeZLqYAC9TYzkuCPiiiSeFz1zy/RgBRKP5o6IBDyoQVvGiigxJ3MKAji4wMNoYExe
/ESd0rCcTLaq5IZo46x1HiJuXRrRmZwqEC8lrWLYkOJhiUezrMfarHzmSn+07NF6p5cO5hSw67v2
LuxachdFcSbJ1ADVyqPMRc++US8EyntCu9CMV9Wd64HvQSoDq0NuMwvSQkyZnbe0lGqg8fOBWqvI
8RraRvsIFyNNH0U16dncah47LTRl7t48ZuFqN2ghrX6KMZ5I6cfBOBM90HiqCzgY+Bk+h08g+8Db
3C+aUSdJ42S33EyQCMzD/WBlLZWMye5+p368PSg6ePRdLo9H4d3QsUye8eNWHvtfNp0BRhCN2bDX
71fLrg8wScHfpgnJvd8uLfwDZqsD8FxuYgE3tl2QoLgPxRpbxuKeLVXmaJeFTDfJZ4O+VNNqTvJu
ACvzyQsrB9vwLxN2QkX3ATgluZBcFuv6G2hLosBUuMp6AweHoStMmLsa8pam9+YHGy9PemmhqEUy
Bvh7zDuhNLUCg6g1yy7PgADkj/xcxgUuk6LI3uhaKA8R8M2u+Fucz+EzfYkp11SCUe29epaVLSd8
ZREDZbWt8t0ssUElgI5Yo4kQ92MVJFyK6Nu4m/hZueFoI0j+NBtNI8rh8jFui9Ex/lSVHDlyf4i3
7VXSt48cAXL/SVRn4g4g5WNGxCiMvdUpSZgbK1p9cRvT2zDP9U07zcfAFNFuni7HaYOpQ5AKMt/t
vfN5F7ILo7QHii/zZb2yC2HhLtsNWEmJmsTJxEGFxUopRuEpfyem7wGOLJ2TpUPF/qUFrBjZHDZ6
Yy66YfVluZg13dXJQVAdjR+/mgesEz/RWs0LBdGaxjAoPA07eOomqYwNdpKqcfcXQSlQrYunGu9R
QGU3aMYsiBkOX/qlrjph75Cvn3HeEW3cyRVprw38rbFDhLEFG5aTL9hLvZZcgAwS39PSq9FYFePC
ptGIWFrq2uLhO23CZiHP3WnO3GM5kFaEwcC6l7rDxppivjyUQhzlIlmMkCULBmbDTDA+dX/xew2U
heg5Rz2O4jl/WDkAkaaKrMLmppXnEbE7tQUoDE6OpsDrvRZnwgbrGQg02FnRFWqdb49rxVNQkoBj
eDlmQjqtqupVoW8WNxmkzZCme7JG2oLxP7Ls+Tk7A9B3y7Y1+Twr1v3UjGaU+ixkX6qChAmvrccD
PLRA2kMR5H+3QvmRkto+/xBLDYGEitpxEx8AVIEy/kdgPQMT05AuiqvBTxG0ZW5fh2o3+cyXfb3v
JruT6dKsHtysxIM8HAW5awPqG82dLunPlx1UJk8KgUuu6qKm2M46GTaBc4GsbvsNknqIHdbCcLeX
Y2cCT2f3+J10iJK+YCg8i//5iEImd/zsJapM/misdtSbxJuAZ6Cd9EB9rRchGJHDvtkoQizXrF09
FThc3RnvmkKnkfBS+2rxuYCRSRTUIoznFTY1wTChfko78Fq1m89MrFZBYf99pcH++MaChMj/78bd
Mo/mB220QA8sPteojIEP7Qg0I+lAMwUHdZPx92zPghaQ7a93NKpuOozri0aJjkFHhhMLdqH53WPS
SZsDKqf3GF/LAgcQoyawUEsQP8235diVsyiL8nkQQAD4c3MQHglZb6B2u7fAtb77NsNJeWh3CmKo
IshihYla8GMdup3V15wspiG7uJBZz3qbRyl3MDnQLr0rSTcVhpoUHAM1clBd2itZg0Xc5HzY994V
BxiyCs9Tj5U7O6EZt2dvG7urjdaJNX0P0hCxRjJ3jxvyQineKwvivXQwwLYnYQS3QldgueLRnr5U
qz92D/mQ6IWBKYpHaN2Gy3xK3FUizTM0W7ZhAjrN6DAvZzt2tkQoBcVvljQKhbRJP6vm8AwpxwzJ
MghtMwkDSHPD5kbdSo7LPyFfuB4luJJkRdk3q9lxZGc+qo29dEg68NxW+99Qxm/0tR+3m/kSfG2A
50WauXagrgCsbQhzXk273SvlaRMwkX6xWCmpPDRCJAQNHyTUj+Xfn/xCaF8G7NRY4sin8FydtuSt
5DEbu5HrXZNf+GyOryLDNAZPfP4o9vngBmGfjH+eeAylqacRXaeUOIyJvZxZvLDTBMv6v+Xt2b66
ywSq7VltwvkY8Z+G7fUrZNRu92YOSUIQQ/c3a39A0HdMsu/3sIbsHkgY0jyXwdszf2Kx8aPP5thW
pEg2SAFsQ/Q8onkaJbHg/CFl+79c0oP0e/2bXwrFDmHQx5j1AmPIC18ghqEUaT6ZZkhJgSaTIRoK
s3AFEp0S72Et/3I9Ob0ffPGeCKHR3iqlIsrPNPlL/oQ37NWGduEsuvUiXHnyfqMN81+eeoG3KDiw
vAuOjrVgbWPQBYbsCragwcv7YxwInTrHQiRHmwvKaiAiXoryWWoLqXCY/rS5osJmI4KjlsPI19uF
/6CGi+5tIhtDfuBupMTdm/iZXHB1KhnJ2SEQESYoAWW4EYag2Ic6HIW71otmhq+3nuyMbyQhkGbs
Bwgtf2JkYlpG7PA2N6vKUWci0/22KT9NwcDzN9RhO8smV9wLWoNpI+bv8SDsY9gcxty7gDXhO2Au
YtQyzQX7skB0ofIwNvl5KuAa7Vwh0ch7hX007Tr41BUCHSqNfZaFxsQi9vGea838RVZbJGkb3KYC
qMsIF/CWGITqQZ1Yx6O7u/QHpGBdSrU2vIlucQ8WsH+ekGujYKM7i/DpEUsH4ZJj6X6ASekY1A0f
sYkHpfGTjr6kKK8rIydlVRALMghQIOldNb+uwDAbeV5/zP9oDQb5tL4dOk2UsSxc8vOS7EEKfJ1s
/9fOg+g/r+TIMVx9kTvJkRPW7h97bpEss33ojpScoAwIk7d+IAAplv59ntrwvhlBV/gzolu07+wn
cgg8w5OKj23SkFBheDVJf8kLKhxWLQBqDbdw0wT1Zz/TzAJQ9OCnkv3mHekLrb1ToMsbqJZVcOwj
UhhXtF0cZ4Zj6FBv4BRUVP15019AJIHQuEJrSUUCLFvCaJpKbBrCMNs4YPrOYWyvL+U6gpKJdm2e
CdYkOYLDwOIkq2k4vVAvXziV/ot9LqpDslUiGnvJZA7DkrBOagTEHWcNaxbmVIZD8YtaMhDgixId
1xMZGBqvBOy/+IHyLCmu0fIprCeOpNUUcy+9wPucVWN4uLKbrA94ehsmdBPKvbwyyxOF2I4A2MxU
O3dtXjFwYy5/IbmujcZ/WQDlCwKymaMqnnUYMW0vx2FwEOYTCB6LHYb0em6nQjwLP/BuuoCEk65d
gA2LsbiYxk7wj6satRSrHsI9MUpHUSUiNwB7mId340VfXjL8XzWrjazMf6MUOqKUzhgfkPX7SyW5
gKY4jGnTFi9xcqirwmdsxkTjiUL/rg5scfi1GBL+AecAzvjE7oitJRiwkvtBjVy1MacAfrJAnDU9
1MktVCQ9XVxJ+HheW8y/usOtsK6HkQSNFwgRyGCkRN/qIfYmtkq6oWa6qOXTROFfK9NcIKGC4wUi
9cV5IbWNKvV/+PG0TQBOOH9xue7pkaT6HKCotHFjGSmUfbP42iab7jZoeNIVkS2laLLA37wWuNos
9iei50KCUMFonNJZVcHmIa4H41hMAc+aggu484fmLho3rpCx3z+JiZNsXZFG0nas5WS2Nl70dbU3
onPM1CGbrrwyuuFGPoY75wTKLZFmOR1lCg3QsHOq9LSSxRSz9dDG5vPcFwrons7c2VseLFEPGSY6
BBAMfvJV3tzNLFgd14u7Obfj3XjGTnwVx2QySfcMjbBVv9D+jBmVYQRldpo/GTbu+sjJbUq++WoD
q1EydFIc/A2dNoytuRbQ+annFFCJcfeL8dhrwytQE1sf4aBTWsRun8xLWFpNstH11rouVE8skY+B
BbEGAIcsg7bQJ2JFu5rQOZb7Ou4DJ1Zd3HzqVUNHmYL/2/kZtYzclDL5TEtjmn4LUUPYSwLZHezI
b8Ih770QK71lweyr5RjbrbXhWHtXCM0KMi1xitFAwCveQ892aJsq7RNIsVdfHTDSsQHN5K9/966g
4tbN7JAz2seDeffIR/RwmSaW/TAbngioEJ8N2g0MHGiZAiXn06rXreTcJUFi5XnZV3pFaPWy9Ubb
ikG3MwmeGdB8HcNil6np6FWgmHE72RAO+8neMLHXgRbWCDsFLzhEf+W6xNRYXzAiXOgO9ByTGc51
IOFPKXVxWXbMthtSE0ZCcg3FixsHCIhjPf35HNjeP8IM5DIc5qeCpapYfcneynxpvsZ+Kj2W3mEO
6wLQGnVubgUrVTjxwj51hnQW2OD4LhpTaaDKw+rTBRUVFNqLy/7dmqnXc9y4IaQDi0cVhnSgXyL8
q6V0dWSSO1Ov56PdMEz52V6+0R+oZEjMxtOXnwOmFeXn7dLZeKOA/oYYQNt7hyC9g3CnpW8882Po
JQOgPfOEG/tRmy1ttkbg/NeqoMRNZ96jKcakbP4UtMDkvn9LLS2qaJj1dzGfXfINb+zPsOep4rnN
PHKSwp/DfhUdkcIGCSpN2yCrsXJFBeq3VTBgkXTV0gl9KmSxhjvIKWUOGTM2f9CUwDYtNksj9cf3
HhsbDwAZfybU+1MZsktm5amNQ4owNo5JqBr/VxlpScA+RRgdJgNcMWB/We8Um2oVdGJvWK/8AAby
E4NaXOk2FE8oHAUDdaaus+IDMeol0reIHgHLTmzO4iOn3/0QthChYqpA+YIUNnmvFlv+iTsDxkwa
wkIkUVLNcN91P2oeIv25lhgHzMqPTmzLmbeFNQEMkHUtQByIvvrjcZ160OISmLge/lW9q8dH/vBo
Mj+87siUvi8CsAeLChmibokz3E1+BAzLOIh562ErOMytMRUyHKMus6pNjDedU5jy/UNci9/m3zvO
ZDA0h4YuGDyjIMozMfnqkwsxBXt+xWICkQ03kztpvOexR0MfBZCs03dLISONFjz9sT7V8XwNP2nI
fbcVoin1HuJ1rI69jGPrPZkPhgsv4jgBM38LyeO0ed3Iu/MLo3zaKujs0CLii7UFlc61MWEoiFHE
Q78wutpOA035Kza5Iv2u683b8zPwrUTmkvW4AvkSZOZTM/7boM9ZWUzDTgHxxkX1rwMi30uBZxAm
DzXjsLKLuVfUjeAk76yzabcUhDS4cBdc3TqNdPD3BkkRZfDeDbtlGplfSdElOoEDw2yItcOWGwf9
YBCZuhQSlH8Z4nRu3m+qD6+bYENIafIwsVK2cdCKbhY863BGcxmAoWOcvsB50P9MCKz6YB30K2hU
2hzmgZUmW15zNmpIvoO3df9rm7OsHulj2lAwBv20VL8Mgf83tdPwZMs2KhSvAo3EGvjYgfwd01a8
V13sbzl3PK73HiR+SL5430ISDrQNrDQTnKweEjDHkw0BZuxsq49xF/8KkS39hUrpzKBgwNkAmtcC
1fq4CR5TqSwk2irZGzAGDXZTUK7ps2/31Vn2YBvEGvjFlYGDVCMsgmAT85uIBecuDF/dHeLEQJ2J
JHlfzHGFEwDVLCT+NBJaoYIQ4jCrUSUCzIR+loaewg3ZlKfYanDlN2camSTt6AmvQYTfTFFU9eJh
ImFWaMGVRMgMgQ++JIxcBs2VPF7g8mL9iE8Tiy980NxHsp0uNNOMrCqccAql13XNsdDev8+ThdW9
d4EO7XZhhSvCNMoOzE9nTq6XWvn8TB7dRCOPUc0ziY2yr4h2OzuczvJy1IFfaXGX9tzHLJYGqqSc
xePfljDt/fYzAc4289cCs/tLo+gwPO0urKhMRn8tyzdDYMeLb5Tk2XSOzcCxdiFaqoR1t6JSPdHh
PGLtGCHgo3p+8tEUy4WJDVm3nLns6nrkg47Jbt6j8pgxTeGxQV8/VVGwORlRY3IVB86nphgEUIdW
IeDORbiwa4zpfEH0LeXsXqEwUmI5PEq+dK4HfBKLuWVo5qvtKIuezKEsoiTWuK7Ai3CUm+a7NKsi
7et1lEY2+GY5UxEkIC+XGMd8V/stTBkjjPlxv3aU3K1D+cIwOnZzJmVfYaHHFgIV2ImO2Sn81vV1
1ft0hok9TwZe9bTwZN+Z7xzROFkuvSIDhn6WSZIm4o4L3ii2KrJkNwFrov/TgJ4bi0E8G4BiDcjZ
0cRkSt02iQeZPguePOdZQrbfE3nA04C2TFBOzmgQVA48NHB5NG9xuH4/X8+Z/BljrXUgbUM1bDgf
2BeFtzfsaDdKhxwHCLnCLqRL5koZ1HymkJUsRBxoIyoFXAVRuVhK9b2PY+oL9U2VuQi9LgqiTv2a
iXYR20eEJea9bgCxfT4JCGdBL+hjYvllH0pqwKLsuSXjvaFpiqeyofMOsosc1vtY2v6OJdJhPHRO
vl4RrP1yF2Q53nto/FBylunDknET8ioJNRKzhC3JgUczVEGhV6KJvac1vPlM6SQ08jcTGDYfM/Bp
EXZTYNbWUlTdX/CG9nGZdIA/2y3gy5tbt5dP/x7u3wPWoKW9ar5JbDc3z1DOlxI3cwQjtXFwer16
iq3MJq3COrOwa6B6wKvCvq8tRfsE4BMvLkgNm2hbyp4scpsz7D8KSJNJyjN7ZYwjRIJYvs+pRkeo
dvwzvGLeWj65VenPfvX/lJjFZCsZc/eZEhGZ8wz5610qXnzpYgjGghrDN1pG7uGP913PL7nPZJN2
y6jKn7Wlat+cA06WreVl3t/1xKa/vwS/sLg9zJp+NtHJds724I9s0tfANNaFez6AYUUzY8FFl/mB
6ubbhSpChHOrk9eyuwr9MYlAa+4unO9PZh5ymXzzqKvrrSXitvCE6e25WIDoGo/pxCg+UqOkva2V
3OlmPkZgRuaekZi90lNtUHWAaTi1tv0tmB4+LN7Q8aIS0YHOQ+hy0lk72Hmg+8vWNWxWJxhTxjne
E3A+39PgeK4wGPp2F5EldCAyxxYSAWyTahZHoP9xjqRGtNIs/AR5TJN5VpQwUl4p/4lSC6SJkwmA
JbPR/G8YxtvtswR/HwHrTPBoPCs7GsMlrisnSK09aH/aaawn0su836o++5Ue2xnuV1kdF1A6UPtP
IsdjnXcYM7R7ISDJFwwaRTEKnkbvOuErsJZejOnVME2lY2yXPLq/0F84uo/zgTQ1xd196+ET9COq
bPldPocXk/dymX4iUw3GKCiT32Ay0yHMbkevN+CNSQr+IgKZojArUiAOgg1NA+XY2RUh4/VOWNwr
2Ejc8doO1WJ9YAR2qbK3T7s4WCkK6Vee8Zfi03NiUBkSOEQqMgpUvfZ/kdxuu9fByjGt8EoFOQKw
l8DKbNYHcYz4Na8jMPaHB9UlY9Ti5qep5S/1Bh+l7OOVWNKN+KA9kCmxwbexA21ZJ1ZHxM9TzUyZ
NpJGRsDkPamKvd4OCqSFBn5zH0kORP8oyUMYRMAmBUro7T2FsmgLbBYMABtvDu5GxpMC2vz/EFoH
yRL6Qf9+Z8n3oZQoc+ZLF0xsTV6ifro2gDhB+ZpJQj3VtmpZkhtfLnn7aOdrdTLngMquiV6TRrqO
LUCthrrTnJK3wviahpP+hLJ3iXcCOZtkfb+pfTl5ChrDEI61rr8u755v329di+soJHWVFJmwYYuT
M2xmwo6ycmgJLu1KCE3x3oYcCAsPEVcE3A/TV2zFoU20KpQEEGXcKQmloE6PIJTmkNRMnENF7uSg
boei0yj0ZOf3obw+lgpgsksrIfZvbA90uk9t0Ms/8VpXHH8oA2t2z9DAJ/5CbdtUoLQdwTpP5FPY
xUn71ZQLvQ+B5DlNJq9jbyYOrLNOcTCeaKFISe753rMXyDJkFo4vK33uXo0odkKNnVZFWn+9pPsp
8vGStG7yOcEF47Lt5LucMubeSP6eJWyL0+CFZMHkBK+ktf0OqybA3LDbvvqJsw8/a2F0x+tn/X/Q
J9qYYZi2jdgCMOm6tOEz208hpMTS5ODhG2Fv8qQV/YGT8kpQhAtOQCBxsbastR07SZMsBOV9h18o
jaJoMpuKRQisGvStPihg+qv2IiQcr1n6+3mViqW+x8TeLSIzAmZbEcVITclXIcfQTgMN/P5ki4iO
Q0lg8YxVxHJ0PIUXxMZtEVDw/xTjE8ofIhTQhYW5fJNsfr+TCxQPz7Lk5eeukqXIFCHaEEBVVjY+
C01925xSDTU2+6aR2O0C1YFyYJutJCfr9aa19YKrp+7ChLO8sCbSpgGqzXbIc0Cr8VguCOeVJWAq
tfj69VdftjR/LnIPKvBS3wawGk6CYvgGhcUVKpyrY4gL22HT521s/e5g5VR9uGB/LAResIqj1xMt
D/twshCzFzQ38jis3BXSxZ0hphJVnpOQICPjZa+bCWDQkLlQ7a4IFA+oEJSzovc4hA4ECcLhcAPm
ATfOswVEg99Om+t854lCUpVOC8NQ+1o9DmCiPIdffKpHiBuj2EAsFGm8A/CkbHpjrAMTpnakOqOS
QH6H5pUa4exI6LTxIVC4l7iLFhlbU0Hs6QWPRMBOyFKSKVIdaaGXeMFeTVYBesA4xQIAQBFOOugV
MjXCYLiLjy/uUwe3r2pT/XJzH5gIyhfBqPPdokeMWPeQ7t4fMqTdt6pnWkMfxbQ0Mw1oW1FZZhME
BNU0urneOKorU7QbH8n6Hg1PWKlKh1lASAQCeComewBlzgjz/YZtmKY1sh422IdDV6dZSJlDNLPT
YteQFfEKkS0zxo8zTOXs1FZBFa/7vtwjf+bUPXbcz4Es5V5mtv8uYQkKKpmztGkR5dhN8socq+CE
WEl8C9x298E648INkw9AMQWmwsSsvnIEAhqDHw1v2p6CWvIRjDt3JHOFbCa7q5lqQOU7HGo7YV/c
VJtW8P9I1D5+/P9gde0LgPO5L4Bgurms7KYLk8FJW82LBEYXe6VZR9atMpmzucgXORdrXOswnyT3
pd+SBjFvdzavs+lbN9G1sCVNYm3/tKutl2T2IPEqogVjLgjN4JEtLnhaDvA0QNjC+FaHy70uDeYI
ps5jlRLeA6PQLf79DX/v/mfrMzOpNlSaa1LTHW4s7Ci55PsbAgOUWWqWkN0QCSM3CbChwJ15tHfq
kSkyOeEvgtFps5B7a/rnKfojpkmN1Ci++VE5Ua9+MbpgZB9RwJCXO3uciSdyEIvmdtKF3nJ8qIF2
J407e7wBOZEhwKPQejhRE9gMaQs/i9x7b9wyXJTvn/qTOoFTrxYOpE8PuKjo0rwZCm4AWiB5fZgH
T2h/qzfyhxvto44AM5QTb2xK75cKTcesXGxTdZwI1BUIyN/ib7xZZFeocusRgnzK8/Ak3Vv3q5ni
PwrworHwfXQ6ldWDaX0v78awXk8xCGR5hLZAPGqerb4AaiD7bpvt3EQFJ7v4ngGSnhtqTWBhk/hT
mZN2ngPzSjeX4tTYRW6iW/HowiRjR/b61uhvMAJw0G3V1ou3WvqdTRgUYQnxGpwjScC8PVL7CZ4E
NLmfO9lYBpwqNFCb7kCOULgQ2dmnAGedkl3DEyjDjjsFkRCbqAbuqNackGZArPV6ftiRy2Cnw9j5
A+A/STaRr8TR0iADTYKGShsRX/jkYBlz+be9lh7r7Iltb0ZWkvjrcr3Cu9+e/hk8g7wc+/41/eZu
Q1+UbcWRdb7kcCEJ5ISa/BbyKGB3MFNM5tYoW6/up8YhYzLPnpntlowZX+wDt2Izin5nsSYP5MeP
MAPmKRjoaoRkrprsuEmAk9rmv1RtrX/Xve44GbZR5iMmhmLBFnqe87thZTT1B+sCd1GVXOxcZa4K
N43YoBS+hYgW3F5LexS/9L89oMF2TOJsVYaHdsGF/mr/3R52a6/EEUk2of+qHA+zMOWHgnGPKB43
9Op9xtODIU2p+Cpj3I7rhyPKsmDiQGCHki2pZMHJ527DQzMNc8EAKH9MpwE3AqtHa2iDywgNfgfy
zGUnjS4wUCKKMahhvf14gIxOzIQPXIaBXINpfNlA+1JUiGgqtsZkWGGGyQ5/10UAPd7qB214B595
mhSlA2UmqnZd1N8UVuDKWcx9nU1LxCyakPzmv4r4NqTaUjhnBtpWsZ5rWKeE7tcgMYl4xcqBUfwK
giAOVA+vlazzFzgw7jIOvGyTfspPKI2ayaRYtidENjOo+1bgQdbsmmLc5hVk/bDPZz/HuLxJBlNo
DQQQ6HLF/hwSKJW4h+ogaGzebj22+MbWGpnJCLkRweRuQOAAvLa+4ObfYTyu45X8NIRgs4Icty7R
NqOzo1L3YLZyFJp8Nm2IHK9KhXhA/7tiSar2f8XdyoqHo4EP8OOCu294ClSVqt15q+7nhlSgFxX+
hgP/M8KgHBx7VZOZKA44qUR/0mbACYCeSLYSh6iz43YsD/6hWneeO5m2OjrH42UrSi5vetgABstN
G+T/F+ec+LCxFx7bHwpFUoroiQInfiBX8Pcic1LbWTfABgdHbCYpsINy7S2Cmgnus4RNY5vUsE5+
27xGwkbSDle7gJWb9+ULq2U8waEzgf8HdNb93J+CGffW0JEHI86P4OQCbR30nuzvqtCBI4zvhbKU
9H5A5xmsCPguI3nC1GEQEwSQsL4PBVaFeZuKimJ8DMgzttnT7MwisB+Lf5OccJsmMYqU1jM12Wtp
ZWvAvYPKhF6wVQwc3i+XRyvGhF7Sj1Rnzi2w9RgKRTJYSoiAKRBrx15jGGUsKr549pOFb0RXcLpj
E3ctj9kXiwdzRgYwd27ULiEu5pyjVvjTk4Vg7cDzoMWvL9Upc2eiJ4s4YmCZxilijn3l7TS8EHTO
oV4I6iX58/w/17P7aPOffjkiLGBtVtZMgAPzwHsE04+xsAvaj1kptoWIZUxoF/WpBEVYBjHtiD2Z
+N9ZLemr5AJjX/uj7sDvNXtjmXyFiqMmrg2/buZonTzmdNU+jH6rHcaC0wK3Tc/3xggz1F/fUINc
8vG1YcCn45fmb9PKF1veXiM9AUX0ytu29zSucuDtzMDem9Ik1HNNctBG3t4/mcSrmmZS+8/wD5wU
a8XSTvCsUDiM6ZjtX4R5M0YoQEc+y6MezPBEdaW1D9gDMYZlZX2jeaKnYOK11/og0y8NvPDX8YKO
7nnBFNhIo1A2ds0WdSrUgqEUH5HD5qpfI2/olLfVbo0yxJBVgRDsiFiuo3wKaCEFPqiAQ7LQY35s
OlQVI4wwQWViNGMVDXpv7WKv3H7MW8AzgBCPa8kT2dW8qMsXio6ENjRpIHxZcVbNt4zWxiwYVDh0
ySTVQMKpHZ441YKkp+3CjGjK8NY8KvTprREpMJgpSMqqGTD4LSBmU4TswOGLky47R0oXmpkcgp+O
q8/a3AMzeRc44Eh482L93B1CP4DNc4NooPthdQf6THYjygqSgXbc/3arTa8LdruE5ZFHd7BskSZu
cn+9YBj5pWrUcISmWMnI3xAmjbJFFuSxBoaBIZDELyF0Dx/zEXliJdIX61E0hrPEiraFpAHwncNH
krVSiFpkF7hpbJrHRkBTr3j9q/lir5m0XKx7rPZ5kcut7bbpvMYEpoCFj8vONb6hzhkoqcTzyf2G
qh9fG+Li3v6h/WA6lbjk+bY0Rxq8nu7j5FpPg4ynqiy/dZ9YZBlcZ6VhfFL7sMCl14L2IPMkH57T
tO/+nZyj9Z5E64fCUYRyuPdSDTzInMOtKFWR/o8NRJJyMpn34BV4avoB9cOT3U4x59qD2TTV2719
zJkvwv6Cg0ejd43grXK3Ek52HBER3r726/4phSLX1/gF+jjcxt+JebH6FvYKTjcUCy4RJbp+R2uV
oDJsOPIKaHrOj1Z42/RmMKdEl7riP1gWt9QreHcYed1qSgtopgtaJwqZjxmWv/HLpvdkVhsJz0Qc
uyV+QHP1e9fuqx5zsxtIJLvv2DvSf8fX69PHGF9qxF4YzxmkvcZGHIfiujM+Jfc6fx3Mb+88c18Z
4ITQcHBIPsQaOWZZw6Wz6hzluOtxjH5kUtIiQeAebel5oGKBfUI3JnImWCvDo6ZFqesxzKMATcHM
81bYBoTWOy50U+evbqITtmHiLFey1cS2mdPBIw3etNzJKpK7l0tZYbeDoCMfHRuF2J955tenzpDi
QQ6X9qRxtnt/88M28xWmofCqgRHj/e5zFCwi+oz2j5I1kYgiaGRXBEpicqkQqaGXZ5UfNnFiTK2Z
2hPMDpxMt84kq0x9OQ9+sBpLD/DWrkSOelYZWGaxBpRNrqWUknNTeJ70lLp02FWrCt8xCas3ZmVI
XOLcEDHF4Man+6oH/nk6n9TqwDPESPJjvvdI8qu5fN5jti1vqQhCW0/jI7ph1u1/yX8PJtcYjM7/
bmsMWmqYcXg+5FN4tkOcCBQUrcViJM0Qrcv0sXsOBJh33/+aaKj5m+lSZTacM4dy+l+Hl2E4Fwvy
4O4uSjVQ03O/EblHp0M0RYx1vhwl8MTvZ5ARmah/VN6uiLkZWNl049bU4OpkRtcyrLeQKvkoQXTQ
CV/wD6HLs8PvTv5++7Iio99AIs1gwyPTRy3IbAc0Hz52akhuEuOTJE2/KnA22OhOsLz/qfzr/h8E
P0VTcdGSE6TAAu9PrIKQImzsQlPvYGVqxaM5WrK9vGzEnKHXI69AWqQNJfD8WlGgEaXxQFcTdQVC
0VjXkkQ3O/L8ZMW333KkRAQhf1lBTJEVChxM0UMD7f5+qJgbxqOK0Ppz+PlJYq0g2C/D9CfotNuT
kaK9ltZdBoxR3o5dvuv5ehtrHz9fOw6F4lt1gnb5VFM5aOEi7/Ja/OQ54WfSIgaqZpR8lsJX0X3O
laydV58yYFf85ivWsTQ+XBoz+bKFDpWNtoWLerN5/aajnhCotWwZQofpFeNm6QMN6A35ja6r66I6
ETLHqFFt+E3RQNeOrjU2lt+GlQrMsH/5DwR2PPKnQQuFgbDF9v87B+wnn4IKtOGD+goLJGzdtLzW
NfPuoDRkPLxDE1Dfnox3NES8TBSu0i4Kk5mjWcizzR1AP3VcNK7wCxCOdYKwh6mDQWgcgNOZ1tQ5
q2QrChNth71jvEJgJEAt8Eaz8PJ6SSqhh8mYEfR2sGwwBI36wGYfs425X9Z7mnCNOU50hM4e19aA
oAiCyA/dDqVXMkKrp1wRTk5p5iyN1iJ9zFEbewv5cj3rjfV2NznKzJkKDFNrQfyhjXO+hZPgJIeg
rjXkZOjXqjMtOZ8tvTpcdWv8JUMIEWbnIPeoj1fZgrh2365JBxAFLeWX7Bn6WfY1JOjXAcEn3VYo
kRd7RD7X6UeGhFOe51YtZZ50PV6GwqW9p7+rSfYy+tIiwHXi/Qkt51gFaAQEsNWt88/G+NEFENMW
+wSqejGf9XoXfr3X+oiBBcoZWlWje4kafR7o3VLB4YohWtKWqvMMLmKOq1qZ0PJ3Ke8cPOOMl+4E
jc0yiVHG9Mvh6bnWzm8y5Drgf5go/84REy6tpwvYROA7tWsAtP+B4C+iPMBvZLQZxFGxAA2/YyLw
DHCtlkYm0WMoM+LltqgQhV3LqgBk5qeoZZvIsmngIPr2U2CdRwm4x2gsMi3n1TxDbK/Eyuk+2rYn
NxS5AuaPEzgYmSOIB3s7E7o0dT/SJ0IovKPbkhbQIB87C0GDcbKckXNzIUpARTErprY1SuM5g+eG
B/3ZzFYLNLSifC3PNd+gQsio0E97ZLvmEswZ7r8xYYRf+H/K7AB8viEfGe7XOo2+TMM34TP8bqH4
53pzINl1cFZ3qVViv8IQiM+i2xbXGaAHH4PWjmIto1G6Sw1inWYvvZ2RrrgkkG2Xve5v9k4/WB0L
uVSMM/LiSrc6QByhf6rkEVtUsZftojvldC5WI0w+NQN05WmUXnukWfFqMm2+cDZLKQDP9BYbnkoR
f+BK8B/s0rqfCmP6Wfs5R7goTvrlIzKOalO+KdVY15WfZsalOx118j4jGl7AItOZMeJv5aUCELoN
6/UlMzRhfsqZlzq7+ZY12ocfI/+iUafGRN9yhSJ4Se6gSd7iMDI+URAXHvIV6X6iWYUfw3pn/V4k
YYngajihHaiMj05bYNCEeLfSFUw73pd0aCDuPdxqNVp2BhkVfco6HlaN5fKFPYRWKtrsYMSCplem
sLenMEvZyEQn5o5r8hYW14evPbAac4PvJDHIV6zIVo1XE/eVW11/b+N6bZVMRObYT+IxR0VHh7zB
jtvIue+ZK6c4rgSMJO1XDBfSqVnBKaB/3UCDagjrhwPswfkHankVaD10LRW7ercxNfIH0oi8lPWk
jOfYeR6xhiNlz/v9LGdnQPnolY8QeC0iRv0Vz0XF5oz5jtY5MsZXI0tl+8LBWokesnisoHK358g+
QtOCGelvRqqZgVi4RRIzx+6nTETiIlRzuE+4klxJHfrRz4DCSTDneO7HmahrxchbR68sAa5eJXAZ
erfcLUyAYlY1zjWJmxMpjaMUvY41YZf/nRnP/JhiDC06qgBPd/CPPgpMD4+OFCfReZoC2ESltbd7
aL0Lg/2asMYD7n+cCPFstKczlnU8inHznEXJVjeL4cyYT6PeyjJqwj/yGilB5ej8sDoYgMrdmcB/
CB6lWEu8bLRgZZ1GHRfuybltYmp6aUkovqxyTVXlCOgwqjkYNcDdDiMb7tpmeonphrZ7wVU7LocN
OXe0+z2vrDbHquJJW4/k4Htp2QmpubA45z1y88qJGs4YQ6ON8A7iR3/1nO0Ols3jldNOHFh7BDYW
gAapt7O7LxhBOFi3/nHXiXL6jjyvEYSHPrCBZDCIutxDpRQ5Aq37+dkiryUkmlGtcDWUS23Qz7QG
eeNvE6QZViSekYObHF7ao53i5Or6qmFLm38n0WMIa51NyjyjBf+IMnyNKpMfw4KCLrtLStlj9kiP
P3v8XqLO+WkmWKmDvi6Ct0TS/1Q7jiEOGUfP+Zx+KSeNZtbOTZ+IVRlkQN8nCcN16O4te71bXP33
jBBEYn4tJ/2JO+FNEJcvB5dJB4iRVfTe8U6sdzbZqOHRqDSDCr0YYtH73+XGS5XRBoBnmQVM2A+i
iziFDfr8p42jRHWoR4u+Y/fBXAl5MhD3iLdYhnljzQ1vebD+CdXJozHEFMV/OacF3a9Rwd5FLTlW
sr/W89GtVWSTIUr2fG/hR4iuAIskwIm7N5Z2EVjNLYYXFV4BGOs8jpmHVDdJicgmSykOQuvLP6dx
MJgUWO/L332Sla+nqrerBgunTCMaZy30vKdPWVXmFyZdL5EaUByCpIZUXvN+qDGZVgcMwraiJXc8
2myTbXLEfAablWvddLk2xEHsbVjxOFCeogbpXhfLLmVjVKMWqGGH1gret3hMAuk10oHMsL0b+IEl
ElapY4cl1vAhmguCaBgz3xIN7BG3acvrh2lW/K4dP7mIh1mxHDm87DDh1grU70ZnS3cjAHTgoIcp
NELgKuRuB6YqNLnVfPBThcvO+unkprT704M4+0uB3BbkUlhti9Oi6UbSbdK+8TeoBu6V93R2xGty
mgen5r2oDC9PUBi3P0os53+yplwPWix0TooAW0MufZ+7Y10u5vEHJiRgG74QU2e/2kC23ZmSyCHO
yPwuXDLENjp3R26S5iTLMefXmT+L7pzBk4G7TLgsdFkgAi8Fr/9QLQgupNVZD0OMDV5IfFShc1kc
1vKBOWIvKsjGjZ3rGE1q+9l26nx0cSj+1a+/kQfmX4LrySg7lEljPm5Tk7WH1UbMlV3vcIIEJAy0
JhupV/EON5j7rOPR3DRUJ04d56jh+Kop8b9xbtHX3Y3X3RBjjrCGz24La8/ZE0K5iHAwoe3nwAHg
LnpqeBuM13KrKsp/9UTVi10e0E6esztBUe6HQQJeei2xnRcsFPCCfMaovuARxlmqEXVFlFsjlevJ
oVjO1qwGsq/mXyKT4viqoH/mzbHCbWq2rSd0qsNeDBcq28EF2IEE6moFTyuA69B7LUZ0Cl8lNIYH
iNwP6ckNzabSRJjAZNo8Ly0rf4j+nEIr9bTFjc5NrUY1TpK2ZYfmL1md7GWXobbhcnguiUKtGUuc
0PJPLk127JRK8ZGFl0HEton5e1eKcSd0VZm+HrsGiuLv7bmB3+1G8DAKC6aTw5EoXVS/26HgDhWo
0+ZDdDnx+2ZeWpLuPiUT+C2GjQfZ5PqgyaTBM8Z7J4qRIHgHdBCxwxEQIV73pD4I2aD2udoScPwX
ArtqTG9EJ28D3WeL+2H4iMojDo84OtbvecTGIIgVtTYA3qi29qgYE4r3/iJBHkQ1sInI1sZIlaP/
eo7sZRJyPPlu+E3s+jgqD8N0sb/aSlWtbdwzsgCalXr9H4x6xQm7QFDsN8eidLYVpAKoVIBOHy5c
wYDNSnAht1igJzcFhMbd5iHbH6lADU6jHp0jtCmbApwFXTXXNFh8eEt1U9QqvTffiwACIjE94e2h
0cn9piffYnonrAngUccTY1nZPKodzrh2y5aekfX8XzKi7XFU+nPI0aYw91uP95k/O2Sh+RqD6MNY
U+G3LtjHMDRDHJic/SxIeFWdtiFjT1mvG7mjyJokT1unmtlsV3VhvslzttKV9xRWfyxc2s6SNNWW
20aGbV9PSKtzeS1b3lWSAMPlKY67c0WF3YqYz0ekq4B+YwfAQvr5HmFZUm/uctZJDXwuG/CqHKxT
3p5o/+VvVXMkJn3ewsDJDeNA8sodbSnLeTva44WAH02lEbBz3970WvFd1md6veb6nwmlFr7pvYIF
2HnVC1Z16hDgtlA558hKzi0es4kjUFEYc3XK6PPZOWyVmTLtHBqih7tfRAa1e353wRPKkLHDCDbK
bimcBCPnjv3mXn+hgW4s31ETvwD+e0Qzat/cHiPuIrpK9GKKaJjeCSHq6gTb/TJVyrNbEU5Ib5m5
SWSnjIhZ0pP6yV8B2imCU6lLwk+G+DQXhy7Fwk8yvmm9wz1jXbiQzGGYYzg4igkhVIyPwsP+72il
tYn12uCPkkHFrVeNJe5scC7oq48OLUCMfGuEyoF7U+U5U47vTf0rCmgNHytXWU8xVYYiZjWzhUgG
H5yL4pnwyagotUDjOVW1B28EZL2iTeHyMuj7iKEPEA9roJIEMPL/uGgqpDapBU5vvcNqFX/RA4vt
9/mWrnpkn3fJwN4JhzJY2Dl02vEh9px2i33rOpomolniePb8ORQm7Gw2kz1MAJOZVFnfbgKEfbqu
NJgt0NiVxJfixMCZRlZML5/eH//zpV8IOaSf/Ftjxq4DekgPd9IGfRt/G6CyHSKFcJ4flvVHLHbf
XNM+kvLpzLB4Fp3ENyRbJ0Cd1TYZnKsgGKPWaw0yR8zZI8NcWO/kuW8tAsyCAzXzQbugJVr/g27P
5wZtK7fnym6nHXt2C+CqUn9hPLfr2aQGhZE1D5uAYFPBi2Gp1qBPNW/nGRZIVJOIMoYcbcZWsPzg
oXQcdJD9SHSmUW8gu1aef2gXAj5VX17vervq2hiKAU+wD0lAtTwK1grFUTq3oTIw9LGc89KXh+I9
AbSGmX0tMzmWAE7e78FSEAK9ENQdMQfTGPxo4aCoPGsr7mnXi9V47SQEox48UVXSAHHfbqPVByu2
mDeXaLVxBllFdMcjeLHLw2rH16t+zZMNmvG6c+G397j2tOPZVrKQkdXvcLcDHt9qha4hgPIwE8yM
sLnsaGQ20iMspfkQGSmyFtVlKxEDQGAV5ueFQcPvK1Gva7TdJ2pkTEbsD7qGmfP3oTBi64hVZMJp
NBAQiYnqEB5MVGuzWBLUmGA3FEN6FvdHGCABE1UTr/go+0UzH60E2ykLS7T1aqutpkzExIW4IfP1
6ZjbMALBArqGJX68+Jb4q6a9eZO684PcjgUDgLqQOCVhq7CJDHGapsq08PQNUSoDqQx6fvebQPLg
ZIHa1fXOZcd1J4SkjNwsJwmhWYuEQDS8wyzGq/sCE+gC9Cjg0oxgriVDuW3l2OWDgONSEUbXnNmG
ZOwppRfQdJzZv/aLRCL/F//e8Ddwa5FDvANlICFlLBlC2fbU9uA4RIYZzrwesvGXLz/03rz3RpnV
v1bSwch20nE0JjYym5OXKYbhL5kBn7NbuNk+b40BVRI/HGoiOMMRMO6v0deG3kWc6FyaJcIfeuCU
yhK9ToBt8L6+q/QVrJLLL0n0IGzE61IjZHkQqXUpoGcB2l9+2MRytHK3RUQBSeyIDBg8HsajXT9e
RCHTFfRCcivv6LRcoqnymxG7pmlyigH3UwIl99RAcrNN7iQDWnqLmnF9VbFs4XVX24yb2rRREyNV
Q0rusBWm7YQVYY60uG8ygUamo0fU0ePBj9zpSo6vfCe2R6gZMzpgNRBqlVARgtDJ54wDJQ48yEna
iu3SCuhgpHqQ8elpx6Z6l6ihtA/nIUE9QE+abCWol2pENBROGPhZ0laAqjh0QMnFXEj7D7xFMC18
F090w32Mvfd4AsvvoekcxYlRqBqm5r/Ai2P1EqutkM0lJzFqiW8zBm0kZyHb0ywap5oeVcj3SGUr
+tz4dyuQ401lhiBu5Qnkaxx4aH1nAwHKzOGVc/zpWWTRqJH+Yd+Q/2C7CMIF11IOVt7e9WQumLtl
/XOEAhlPRP7tC2O2iQJfuDoZ4++gx516uJxkytz3PZINy6jD6nFtsFzAhjebrQ1efycUg1IVueMS
avVlhdRVfJ5zzZU6jpsz+4hwW55w32cDuNMe+ukRg0/hZSledn95SkL1oStCU+s78VEcxijVVSAC
NEmf1sKHeXlQ39MacNyfHY3/s1F5ppE2X/CrXolmSYxcK2jxtmXxiZJjEgYeOtifpRM/yFZphAAK
IEsogqA9ZJiL7xHPHHR7DvXap6sHDpm6sbCgLIBVux+36prY+MXuPdP8PdOSItv8FQauPKfiglMm
pnNAy0vj4a+431WwL7jj8SPiaYxMVatIsXl9JOMC0jRAzdfJuhFm1EO9jDlvhI/7zEJZz1dD2dK/
Nwd541EXUzVlpx2+Ja+KHXBg7HW1fweyX8sXVnzFxrBoCx88ScgWejIocBiG2BgCLDD5usgaX96M
NBWYdmJgRvVPzbr3LfLZZ1BsDNT1KSgaNRgb4AoncBGQfLBIQRLLC3cskW8uKLi4fT6txQhv9JFD
7sxVA43pBX2nOxM26Bduz9h15tXXoWzzUhXtP5K5vNuBmgSIy5Qh0zCUbdk3jhsf5dyjsIydvnyA
lYdn2WBuZuPlm+gv3KJ0jY0YKXJHRmnJkRVxIpnw/JXihXx6w0ln0VDjER9NEXA5FjykZ2Kx5xUx
WgmAQ7zRr3DvPgD0EXLXRMQqk6cHDWPjaGDGDbiT9gQnb/Nqlslcnpp5CQzHMmB4P6HHQzBo68Hx
tIG1CWMJi/evOQt/uzMS18e+4U064QZnoKTJdpp6xmb407QjW41F/kKi4+w5+VQUeI71dJtYLN9/
+y64MVbfoY45QKIaiWwbJvpmwPYkekD1N4D/Iu0tN4tYsrApOBOvkzHXJGA7ySqZeMZxBt9KWiCH
P52/Za5XeDXXnHEoVPqI+JfjVH+b7me89bOfOOupjGcqXa21gHET9U9hDMTpDI1TU8r3SLiUgR2Y
5/iHSxbV0/5NLS+oSpxnRuRvXHSUF8GjRikfkXwEk4j+uWmwSIPZ47yQuEtzDQ2OdXZoO16q+WkO
LXjeFk01et5zD8LU48Vp+W+J/zN3Ck/xF3+xFoattAezE/fiCy/c/wZbWMAdrb5c3N/wMvLXg+30
xe/9OO8YdoDhkR9ULVFBbS8aQ+rIHLl02W2J6TDVo6TkPGUkIkQtRugeEhZYVyC8XcDS8n8ps+sf
DxwpbE1l8KQFwLHH1nuBRk1CiGpt1NhYwboKmcKOQ49pTwk9jeManKm5fwJehfaKogqI3wLAVjON
8kFrrVzcMNog0htFsqH6WPhnkp4uEDAggGz2nWDCDlIeMlW8csT1EoCzycm2TbxvavRVIWcrxwkq
osQx77D+PIma+FcZnxvUBIa5uORFXYR44liMISBbJEF+5XK8RPhw1utLOVyzOYzdFS0FSbXOA4cx
AQEdzsIGKmxpF7LJ2CdYt6Yl1HKMsXfVtUTRRtD+s2Gd0cylVlmLDOeFOZNEH5SGedblWuqf6MdR
Bajf1q8ktPG0Z6ZJsGosFj46N27WF3V2BTWaREupUw+mzrvtM2QqbQ/4ydBVi7SeiZK866aUv5uO
VcPF6NHCrsalIYqfgKqb8IvMeBzhAMo2fGST0sm8Y3Pe3q50WTsXPXpnx91gS4nht/FNt+8r/gHW
IKRqPL2S1ei2QyaU0TABNTbBPe5l3Zzy4MtESH6ZYoVdtYVCI8f7Wg4/hr+fbJvcDNgCABdlUC2i
Z/oasK9kq7DfP61t4AXIWrjdr3Q9lguXLb5b9l9x2w5lRmKTiTFqQO3NWGsVPa/wT843DXJ83c0D
Y/vVUphwxKbzPOLVz3c6rB2/u6tK84cS+/bZQKGbCxMp+afCE1UNNjNXU+N2nK9srNi2g0j1lctu
nA8GnPZhNTxvJgjKFw+SDgM3SFjNIXAOjCN7BjYzhBWrIkFi51tHX5RLx1HBW/CYHGknmi2eb351
wU1XpNhTr0Fd58Wnl/303uLN38N8b8ppmkyqzuXZuhnpxLutXd4mskDaCuVrhmuIBaRjZ3XsFgth
1cJcIPv7Wz7XUoShYhENW5VHf7s4DtMC0t64vCjniuL9b2Vglf6O6CeamJkYGTkn4ooQk7/dnxUz
FC2a5OiATHukoUqbCaFInwIruL1NMzWE40/irYTf4DmCkmzlBeZLMI7MPFsxu0RKKDK/a4LYIfPh
kJ8TLe854aEWahKp+dzHgNGMvwHabi9U4kdy4eoDD3ncK6QUpW4N0j73s40JaXcC5+gIGkW5rpms
kawATcEUMdcEb/iJ7d8Ptg3sMi22KXNwYZeSdIyz0n3hYWjNlsAHg/aWB7pJ3ONNAV9FdeOjkY0i
HDJuD8U+RLNOk2ftzrPG2EX2cECliz1N8tVMd7tv06Flu/mDmRz/dXY9nINPjcyG2+FrJn8X3X6Z
aLU+PjThOdnuahEuuiz/wR0J9f6ms8Yz7PiGK0DYPQ9+goi/sQGO2U8I/GYYRvSSK7Nct8wC7XKX
Sse8IeFJRpbF7SIazFeNnp5PNSpTgrhy/sBua51xUEDoW1bnXRqKnJWjtvTUV9nvwnskEYiPRIUX
t4Ugo8dncRLch5nKzoFWFPA12sQzy2/DQGNnMWqXJMPWv++Hr7yuJz2EoTREdTNtDwndkPVGrvHN
aNwiUULsQR0wjVcuz+nBvTRJ/rowEQjdGEClBLz4vEh6MREUMn1pjo64ZzDwxNN85K3CbMgcvEi9
APPF6M+FnIUMTkH6epM+Q9rE74q3DMLRfh6fu8wpjfWxivwwwC76xX1z033FP1M0mbK+vStbH37T
v5zfle6wpMaNasT60GnrbVOBhrEF1T+5Z5YeXrfhXY9RbEFkdL+oReivfpdJUat5KUG3WrEqJ+9X
CiLOgUbfa4Ovvj7E83Dh6sG+SRjTcj3q6Y4plPiN4xpwgjF87VDc09o8sYeZbzJs2K68fJRHaQm8
cdxbZBCOl6DPRckDbf7bHPIoLrwdOHFubcYMxhYCkjKAHNBK0lM/+uEWuELN4GvkJYyjN7hOb8TQ
5F/pIETFcmOLaFlHnBhwPhM4px5wUL6hyBPdRZEimzgyLjX3RY0FvXcfyqAoVUbAcDzVargSR1Cf
WJcPPm1KVJpPbP6cR7PQlNRW93gfhgFaFEtKeBtDoAgWb5+pZCMlTgpEUZdfWjN/GGDjCWfT7NH5
tMD2tYjib2JtH09VGIW2Ho6Vqsuy4iHgXI3qF/AaB3R03v0WKIimA8nmgnjILln21JzxKwUKnOEC
iIDAPyrnBwqS7u7kiLt7GCw0wu0Qk1fzBzRS3Stjocnku7uNLypFxt1jqSfsYaM5MqR9N5ivu+YK
M6hC1e6LV3vnVn0ipHYM1Al/4msD1h4EupM536aEpCXwg9OlrVvG3eEFjI4zgQQVicRmdTDHzCZZ
qvw0iKNVwkqzFx5w8cgB+xPx62b4Pc7py65s/umLVMAH084eMqY5pN8d710kjHA0JwoVbh5qzt3Z
+C2/nNzKvdg9MO6uy7pM39wmPrmjJmvn9JvGQDTf3/yZgG+iJErqPEowcZ4v8+54kODmNDDJTR8a
TIjAX/fCGNZnsgcaz1Z4x29MVksJKJit9xu8Vzzvb9pr1PTLxwwFDarJpCzC9Q6QDLRLo0D1pyiU
7zybXxC3Psw84aAgazqjN8lsRvrA39jACUjBI1Asb1DI6KhSbyEucBDCl1wh4jxQu127DBIr/ACg
JhKUim0QVjbQX0DWdKtho1BiygP9WT21RVsVs6kDniXl7JLhiL7q67mfbL01e+kfpZ/L4NAsAMSo
MwTJSqUiFMN5FgIo8RjgGE6/S71sEJM8P3gglwzaqfyJRtXcIndwMyxokc7rJpkU0lhCftFBrBcq
Sw8mlgClpMcUd3b3A7Lw9ijgzI04KKZiygHRoK400lhxhNg0OEb+kPPxXhift+fcvVrN/JMPuGxI
pRhIceQcvnZOq4yB0R41Cqyj3jhFsN8d2Sk8eue0wCGYS0dVQDjHi/O/L8fdhOJHtceIqK5rE/rE
cYi278/3HMnbnLuUbIJ6tt6vXDyH/RxNsb8i2VYMOkp9frcLf3I831pMfeb8R4rfyV+03MjZUrUF
pW6bmtP+12DsF/FVlBnlaBYQEmFlFlsVhEKu97QqfqxxGvgZ6XI4XbcqrE3wQ8GnFv8ySOjC6f0D
4lbDhP5NFrUCjcBIcH9H3I3NW0HUVlXvCDF85nvNuCYtBNxlaTqGHLmlYH4i1JCQHUNBBFni/Tam
L1UFJny5oClygUtW2gjzQOtKmvQaDtLzJoz7CjkY7FuVOp1t0sVBenTGEqssTniqzUtVyAd6bn76
eAytfest8dtcunMY83cB0rDM1UQtewSq426UZsx8gwgLsWl7P+xMfR/hxpPUJX53f4JakhZ+3D9O
DPIPllnAACAYf4LvXH60BqMEXg0HtuFk/2+lO+hEnCHwbTw/btP3AxeBXoxW6jMX3xOqcM59u99J
+dbWbdcpF2dy4iDxTsRcSE4OvXN3CcKA+54cISRi6LQflyjKeeVYTon27TeoLRPUE3784FPl1jfv
eWa0kegha2SBQ4M8V8KW1ibWV0sAqRE8yI3XI96t4DgdxUzDIFxHLtnH/j822nV46Vmw64KnaD5j
JINupICkK8/bIfjtJ+qUvuiEIq4xe6Olh34TUMOWdgPjGQElUyXjNn69Y/4jEuiiI/cCwwmARJak
4IZwCqUZLvSah3WV9SNGah42WFsqDr40I6MHK2M/fB3SRjxUqu+JRM9/mmkef+mW2uiBpIrs71N1
BQ2u/E94rJhbL1Gk9doMMgPeASyNUW5ezyAOZzMX+OdimP8i+IuUqQyXoaDzsUTw0DlVWbVRe0Fk
6y0O8gWFHrWzCKiSlVGeD7AaymRPBLXtlCoP1ZoZaFCPhgF6X8OXroVWanlRBIMLs9HqmMTqUnWJ
Zd8RFqvbgpKdccWaLAsmz93FcSk4coK6AXp0A/Nx57mPXYg34YudA3DHVPDVhtF2wxzGDq0eHlSm
1ZWq/SEOHdrIyKebNgfAaf39MeQMLDZUr+4NxWlFITZdkhULgn07nbD5SLqt4BKg6p6Wg4JE9Upr
CSZqw5tBdH+FibjMcmg0awjorazzaoOLoJ0nQvjAxhDKbNv9UQhcHfn6p1DklaDPTmthxFS+FIQx
+C7PCkwixYupN9eaQ77hxdJoGv/CRME4h6ZlbqtIe2+gRjbDtOGD+8PUyQus+F2DCJwKBztTSLDY
SLVCtsZlY/l1CFHYMLtPyp4XeVQ079Yol41PWf/YbOieL0MXJ9yB3JUWtZOgv693DMLvAbK7BXaM
f/TmyIV2iSNReBKLWnPSSAUA9utrrbOTgaODsekAQV9jH9LKEL7ErIk3VKS6iJuH9HZrf4/DekyE
ZxyK7cXVnJwylcC9DSVRISuiS+3UncgldpXxx1qMg4r4oZrveu/L71z3plMYaW/EzD+xYcSnvjEB
Xg4+XMowibAlFAgPDZJ/aeEjiDT+i6OgjRC6lIzg0hYJTO5g6qUuD7i+W7zQSoN1TB/kqkQU+oza
aEA3aiNzRMopqHzBeYiRxsL5+1RihQ7ZLyfMiWbpEko93rRx4n/djWb4mWs4EoCg2vn/3LG8XZ4N
IsIAOHRxbBov+E6IKzfcuxfaU5Ns2TH3KZUAOngRDMUrgKLwxdQgtbZ3nRTU8+SESOSlXLiiSLce
MIKcCAURnalfGhHFhYG/thohxpzOimRGtF3uhhiZ2OadoW9iWduYuMPmGXTJa4oxfcmwLrG4pTZ/
17dg0bCVN0FKpyHg6mNzaSnlwEBvH83D8052pGAp13sYPPSzBo4KCbyvWcaM4UnJdzJWQ6qONMX+
F6JAzNvZn7ByIGpfepCbKTiH9Nj36NO+2qUYj90U6rVgeQrLt5NbZ/jwFW3MGgalKWGIlvxhEfho
z3x+a2wBiwkqURe/4OdeDK4TuapjDG8BeluDvRbJDedpLt2Nm5VG+mjHOLM+mSLihsHExLR7gIYq
LTPTVQrySsVxkZn6FPp1aC1XsUEH7xoy1n1Rmed/Jl3N7dJ9TYBh4B1QW4oG9adPiL2FWDRwy3E2
bgr0BH+bFhnSvsG4YSMtW8VIqgu0apqk4Jt6ABAEwGxFM5c15caxlB8Q7zilv8qku4IqqZi8KWld
bSo7Dtk/M9h9cppPaYzQlPQrI9F3yZnY3AXDB9IX0ljR22nOzP8t5faCBNrRhlVGm+DurFbc9lcp
1ZZ3ufk4VRPMjtaonnjFKIjH+JGY6o9Ou6haLLEvs9iKZX02g1PJRdLEpdzEUW+gsQ7rSK4b/lMA
1dCgmVMU8A6xhY+0LEgYEwTjA39hPUvLJdTdppUT9NJsAM0P8Ef7j64WPUhj1y68x+g9u3RHUbVA
KN64AgHUrKvP9qAgJb5ylrV5QfksqqCbMv35Q/zVJmwl1Jauu65Hi//yIukoE7PQiUV21ZgnXqJx
34fsIr66lSVsQC7rwtkvFZW8i16VFepXBsD1Hbns4ZH1dUeIHu3MUTyzsLuijsK4KIb7SdLHDFb1
B/zDHbC8UMwbO9S8W+qFDfrzZUFkN1SBGpaRRWlar5Ef7Fegew8FnKTHlK99zTHdZcR98ClUeUWT
sKoxmZqo439UYFBJOqvCoWR2/iWAzt4LxTs1sF8zen486DNdtT7U2THUbkxTAdkvY60LXiGZmE+a
hQ3e39lOeKbawUQ7f2TRsqNY2+xfIzWIwnEVxwblWx5ZTlv2p00tbzdf39KHstUcbY3EWbMJbyO/
CyjcQezv00Zka6md4jWx+dI9fMUSedhQSTXAA4KRVujlulpd9xgKObMJ2p0jBOZcE9VAFE84EevJ
sX27wjnlgn0eQmqloTwCIU6swyyxjE8Rpn1HMbWlGIKCAnRUjqU6s75OJsdjZs8irCP5s7OwytsB
njCflcCe0w9cjZAGi3j0tjeAb1iFQRn3KNRw5nrcdobMWdOfeMZjnqa6pkM/l7JIfLCRUxifRIDv
pEsZ595mZqE3NjqvNM3bpZBfPJdnErVCkk8WANT3TTGQLixhBnKSQVVOps4oB68+iAFopb3aB2XV
FcFzJWoD/JYWMbwsiAjaMP0G3ElhTWSVAp357FWz9Sl5S7hWdj+yA9G0koKpy7mmA9y/+2qPEjAq
PoTuCu/A4fsIwmsw182052HegSTtrnwdynmvvg4kAB4mdKEJ6yqdD2gfM5lU1W7MrJojx04oosEe
hXalLAqOm8vFmXw1WBKwaLi77JkyCxScEa2mbliqW10TgFNZ5TEYC1GFBsrOnyknsOQ0Rw3V31Md
DEYxj6fU97po7ZUay+k4uxsKrYp8/jjo36COyyyBYQxeFo/AvXlv6rPR6TM4VIoqFGsjUmEjzKn9
h95JJQdhpx8DMfmZ9hc6qBkw9psHcKJLq7NCs1oR317HBLCf1gaCWxj+307d0w2R72JmrWj861CE
uDOa+WZZ6drGIiW4mdEmknUlZ1YDKpbSJzZfm12CH/J8cA2UUIOfTZ6dpDK84q/A0VZ6U6/WygFh
f+tD0pKmek4qQGHufkY5c0ClI3Gg24hNxJKvXi10OmFFwjRwqYzpIf29upyIRL2ZYWJSxLSpfY/9
j0bXILcfOAQjiVqGo2H0IALh2OsSsCogsntjc+Qgr2xrTp0SYMnqb/QmQ71G43r+XOzNy3ua7S5O
yiCOAMGXktVVrZMoxRXBguL97UaxsKqEiPdbUCSU8YW+Jk4NdkYSxRZuvemzmmRHRlmC9RNygdNj
WXOFj9XN1NrimZb0JAHvb0Lqo4+tfrBHGfCvvkyJ4q4T2rajIc9Kr9vU4h4r9JdS4oaSwrbOhP8i
uMpIZQveSgUXdKCTDdxKdpaUL6YTcyRTAgGw1T93yzNvSFBrNNIRconY4aPMlrLvNXmFAdQyjn4S
uIOtY7+Z3I3vFimoQ6SqLu8EINtfxpUMzIxqXt6xsS0gyuT+00/sFLYZ5Ic6nq6Bd0h/0XtDIlIX
FcOiuH9WDKa1PhDiqYPz0tW5JlQTvZCoapF1GqgAVu85n1b1iBsjfmI+nIRncI2sncP4GmRGQ6AK
LMwS2U+OW2DORRmLLOWOlZtmHbz49hui1r4fYwJQEl86024M2HK7e75uXGRv0xVR7zSCXGvAr9IP
sFfUzqkR2b7NRlvW5m5kAJ4SM4KbL5gE59EX1ko1ygJjUxLamE0Kybd9jk7zRo0b93MeT2uynQTz
ZLKvQL7wHZs8dPo0dkhKeTMQjqf9Qx8kToE0U5pPgVlaeSx5LT1EQ7eRMedjzGxmrOEOF/Hn0gGx
v0qrJp8eeS6zUkSqAKTWrwjGmM6s4EAWb1yolefs3FheFgeieZXP1kinn3+kQhHy37pJ/cNg+9KD
bLSArDzFZXpKNtNvzLpWVjtp9eyq+AZP51OPex2p7JlqLvzViHp4rOq0dh/R/ZvYRTsgxu7bSqY4
HdoqcJFJwT9q8+aRnIdADZYFNGNKTFw09BVM23ilTiiGO3IvGXCl9PWmw9MBqy1/Q/GBcczl1gOb
4D0eumCaA45Ya5dwfB1yNNjRC0cOGcc0cBf5h1XtJhNCgDXbZ8oE5KDVP86uJD6Hu9soUXmTt1ve
6UEsyrxNZMz8qkIl5m/UOiiG6nnD1mjtNAUI5KdX2iZkYwoowFcvYmZy2DKCQhxqFr4xomJCwzwE
B/UiXlNZIcomHUNsJYwJYNIqsv9L1qVjssQpRjBRpj1OGVHfi31VUaSi/APNu+ZFDNpot/i2krxf
1p3SyrB67ysEL6dTKSKkgbArJ2furEb7+cCRsQdcMuK7ODb4FOmqDLHmhsNIaM646CZBMPV5oviI
UyyqvsjFjn6dDutSCcUq/nxzNLb1RhSFj69RmD+sK4sYtBchgpiyoXIU22CMzubWp2dxZzumj6Oy
dODaU3OAyHFXCsBSZp5+vQ+jyhGEzXfHqxJfwN/BPGwE61c+qmfQOi6s1p+qM6EJx//wC9gPiMlt
ET4UnjFSZWR2T6c4qIIIRKZKGr4EHponf0xg7lLuSEQ+7eg1oNa26X13qjIStKaaxBo1y4L+Uujw
cQllqM8vUygXeuuqFUPdVJFCBw7BxIFTsuP9amamWrQIKQVjb7i09jkA40vHirzN7rpd92kbwdnL
P6b5mPodLqgAQDjfJEeSxibISjsB/LnYYeia6Lo0Flkywy31Ka8oFJYBOqQkw/xeRceWtLAwJFgM
EL2RfCvDGGX35frZol17YThBJSkh2fKq2HIShzJuUr69Ht3FZuxphuLNao3O+BdfXlmhoEVxQ3Fy
lkYE35J5J8paPK13U4GXMWSWvV2s4R75gltRW3v4uqGoWXeQ0k42Cpgbjzv22UyYYX2aqe2FHgWb
Axo48RDHszmOc9ineEasazEym19GethxCWHbtuBuuhhxUuo+UQZnaHCmhhlKoYeEeQG2IOFvjOsZ
qRFglNH2imhzSYERXwaBbFdNkCTYHzwGhN4sE4O+RrE+wdNM5z3LzQqeDSqqebu2E3Raqbpx/tMF
hjZICyXiDNN1ngKbBPggkqCeVpEO2b3+JXOolvjZXPqZ0pJnmSRXIsnIlfd2emr2zXMIIGA/F90W
MyakUNvl5Z0m9Qp2VcouAwKNuc5I1psIYwVjDWh8zxwC0PzxpJuDPG1kkt97mYxA6GXH05vtLN6x
gRaX8Abio+uLDvJYHGPhBDdzrfpn1AHTV+SJiU/ze9vAiKzd1QCNvNe/7CzC1swvwqETdfb+GiTC
BQZyGEetMUtPS6Q3Lab7/rSwQ12M24Q+grLf5PVJCKfQ4P0MhPMZzWyLFSES0pWipAgBSZs0+nKq
jjoa+2UABWFN+P5+/QJlhaXMjsi9C0PphrNQizZ9gvl4ycOO3cEoRpkrLjHT+Gcav5H9iHgozEYO
9G2tRBLKUJAybGINVrooX7gBnmrJKzjWXZbKHHpUeo6GbtI4XQ/z9n3TAqRvjkGWr0UVlf4/RP5t
nUvzO7nrqXy6eE78RXVtuKos8ESlb3X4fv75phyRMFOMZWMaWSt3nAx3731BtGENA3+mross0bp9
lEN1Wae+b9VrKlbev5T9RhCY4QVe/mXg0cAxzMXABn22wB7ltFwslLfJnG2uEXw1yyktGheC9WZ+
8Jly+o0OnEkciU0k5KgfVXiYTfMpSWPtPPjijdI3sKVdnbsgLGUXatmN/aYLVFqzhJgwZvKQ3rRM
Dr1Y9rMNy5P3p6V+KQxIUJ6+1eKVXChX8EUrAtkMRzJkjE9YhEs9B4/pelgYHashZAH71h0eIkwH
+NH5epfod8udBDZp6gJ2l9MPsktFwGoF5q5tmvAUqvdh8/6boA7g7J0zeBlW9Bk9sOSPlzbqj3ke
6+BBVPTabpFWb0dRd3j2KA8fSQLIvO2RZ7IFOaWORzJuwRYUlF2t872LxRFOh5zSchOR/juEDhc/
Gv8Ey3h96977lfZVV8ixr2SkJTYUIBA7IGABhTsP5t5mxMWOKl6nG+kjEm4Rd9S5rEbbs1OxuLBR
7pF9eZAKapFvnGdmAD7xCP74EuOztWRONg4bsrzI2GlsLma/RMNcpBgRSNKAR08U98CGgt64RFUU
eC1f+huc880pzaKc6f/PniWk7EERLtNwL2tJ7J5Xdi1yiQvV8v6xeeOH4XRosvYmSDSYa4yk6V5w
GQycOO5Pl9R6a86EGuerdOJvrLNYJfDGdDo2DKswdDH9LkPKsBLA1xkapdnVk9ogvTVryEGsHtRA
dQoupGfYw/B73l2buKW2KqA4kgfZRad/aal7n8YGrvPqznR3QoJm0FuonWHCpSRckCpJuzCYmpv7
ZIZZppUvxEGXDgd/DfESeUqUatuKqtUBEpgP8SukIk2DdayPAKLlqCZHIYYmObVLgXRq5Sv0YTCJ
HIhTdxD7FuikcsWOftoWRpjCCq0R5CwBdd2I8vFYHE2iohGpktNjFRlGnOaRd0e8R8HTc6Qjo+ax
hFNAMsOxHNdUpgK38h+pWaPxowiAwfo9ccHuWfkFH9ToBVbttfZU8Ua5oM2bqquJb0nt2T5M9S6B
pvXEz1PsweTncBw7ox9T/CwQ6F5adbzLxpLILj5628F+t6QDBhciqe0DIs/yLR9B+IlJ8BGRXCEe
L5+KRBdJk7Rb5dMbKjAFVgHolM1ak/N4xnrWpDOn6M9tnjlPeh1WjdvsQaS/xesi589eUcPctTSp
NMyKfduOFHoLzrLlZ6YPqmMZrLnM8wbXEcLLdJtZaojnm55kxIGP0CPK46apEygAi9IirPSRVuYe
ni939Y9sKNO5qNmXtpUkUFfceFlOEAO5+nJSoiWYEkhRg+6k8dHwYr3DrvPFKHJNqt80jSSxodrp
Gv/02Z1uRtBGTC+sHpBnG1nJpMvXVALnlMya3/Bpp9enQG1iUJ56xm9UYhjkMqbWPZvvDf1OVK0t
uUI50d0qkJMqgaJQltGriZmbdR5vAwSfUKCBQGeCqwb9FuGH5lecq4nLBRTxNNAHe406Zoth6L4q
LR+w7qGmsHKO99BtErF2eBctLqN4wuPcA2U7+cjhm8uc7MZ2CbBSC4NIiTOGPGCg0OcDehNTPbCL
ftwt8MZMfNE5B4B2ss1ykHqiVkWzajoj41kavmPMaPXHeWD8L7+ErYL5xDgvVvk8Pr1M9vabYd5/
+VKSysp9UwVRUH3xef+14iQQlqTwYgRlRIIDo8t90cje4QyoJkMynzdx/nWEm2e2tNe4qSbtCjuI
SZN2SDP+iJ50eWlYpgS2BAMpLOAeoB3kSPR6f6eB+QyCKiGr1J0dseT7aEiT/Pco9IP+d1AfJGy4
78za5bQbUMIt/0PBBoRzfy0f5RKAghggJ2F1nOKZ4aOzVtOyKmE3gLMEg77hFhWxSnzntKvU9ttl
RovupcNkez/gnCdIufgWUapUDYUPZz+XctLobFvha0uIpQp6GaDH4opvPhBF5gUf0jwR/38cGjSu
Q152LQHFayLsdo6ogr8dQyZayJl2eH40zjn14gryposYgSb70s+5S2HmvlX+oCQwzNONC5VA20DZ
td4GAtprz1X4akOVZq/YHYcewAFfJbn3SD9Fr0BUPKOW66qqN9NPUfnBsyB7TQ/+dWQImxkeWQ+l
/x3o2ntE1UXeE9VBlRBm2kWVQ8yy0JfMwe2Y6oh1BLb1QyQQxGDaQhR53dpTz/Wc3kzZGN4wVW+L
5teYnbF4HxB+FIGaz5dAOeUO5HVyhKQC3DJHcHfyzK/RTdOYOnFSGRQHlKtXGmznkvBS8z+Xj0gO
LK2OwgtThJSeQQS0MrUZ245fw/fXO7UcqHPbriFZ/g6aU9J9UW5AsshUPSkWpdRgCfjCRZYYsNLP
TvHZBY2EUpEooYM9bup1QISDlmWmzrvGWWIyCnWsahA9G8ACn+ypXsyuvC/2cGIas32fkvJGqVjw
+Fdtcxe9YgkQwKbTiY0Djj6xHNxlZVyuJFq4v5MzS1bsedy2IuDATBpGC0uEHn7uwxVmIm6dCf/y
c4Ar6t/5p0B9Ps8YJd1zPgg7WdYIQuNGlgudIMuHVcGVF//UwM7qyerSuVcBK7OZpiAamP4+7WeW
kwIJRVUeWbesAD5eOP++RyEnGV1Pg8XWtqM4Wn5yg0c6mPYWkCGrYcFjs/ixx/VsCI3HR2/hU34N
zdlxMIi33equJqfdXg/7BDoxINzQ4V0rX7Rd0ikkRcKm2K1wAMwQiVah1k11QgaxVP8YHsfJPY9v
DA+o035SRZ7JdcDDawK6vCbqhZN15ifXwtAhm+vHQD7In+cal6kd7nmtRxyKuikT4tu+Cj4ELnAV
/LExEd6+m/oiYY7lrLBcH89FMPayBOnK7geZey55lrQ5gsU3meVEVJxH02JZ6zfcmifdNfDCIC4E
WCgyUEbfzQCewnYb/pAIJnbTRQGb0djmLBwN/v23u8MtwvOEKEB4CRmjQwD/OAfU2U4sXUn70/tE
myhKTTRkKITHFytcUOITvD9VefELZcsBfPYf4qvEqCyEuHzK/kO9o+O5BMaN3veQ1eh10l6zweBQ
G9n2wrJUOaotytOHFYSvT/PLwTYr0ZrAirIF/QOmuKW72dOL4eYegOuYRiStjAjLbHJTGqZ0toZX
mC24y0LEV1h3I3N7OzSfWEesCYB1GPoeVIH67rqnaZ3n/uY65sxSDdUy8y4maW0QzSf7+8i4pfk0
KmfMbaK1y0w8cyFDeO+VbztcU/N3djLH4uxR+1gNrjiuTGfi7wNLozpQOvxsz4SBHG94VmAFYV2W
dLlaq8gOlOQptSWLKBKtkQpCe86TWs9CBZUgrYhYaL0STQzfMPLNxFfybOgKuOxm1CKI8bw58nCO
iVghITAq19/H0MyW4yFGzCEFmGhvOodosZBc16YyYqkffKlDcP7BAGO3wzFlvaQtNZ3jeWwMd8Fk
Y/I+ibJHBtBew2IGFGolsuNWrxjpgEcqaryRLUmlgVKLXat5jE98lGCLa49HJzGzYFyDN0XHOgzE
zjsSPz2tyEQ3h3P1TnY+nqv36hH81x+RLtnIeZzeuT6HptEXBaXTHTTaTLStCdKEriZnH7BhFess
J49vRExq8uO0P2YAcRcSzP9svgwEKaZMZ94+QEqBOn5UvfjFl9B5TVIbUN2ruoxxkeUwjjoMzcU5
2Xt9tMfUssUEpQsXfzPjrxxHWjQf4kAyPe2qI51LvZrTpooY2Wbdm5lLEf2FBo3GmjwympmRAcJV
Xq/TX+Hx6vmZltZCGg15f/CVdTOqbBVYZno+FbUMS+qms4eYnLhcbWWnzmH80M7TleWLV4XhMPXI
L1oxnNzSehJG5jJW+z0B+2hPgHj60uX3F/2R5mLVrNpBrCNRahYx83qciL9XQvC94sFITcv5O5JG
FBPtXjWnBLRbZbUUgggzfS5oy/qHmHtxXWKEVKUw6/mgyW4ySELvVqbqYo8pX0LucLP4y3U6uBOZ
JgElQxPhjkdASmYE/+fpZgzGUfXSAqW2nbcpBxu6pSZn1oz5iyqaAKKGiluAEqGWgGD8P7MoneLI
dW4/Rtg0kdxoybt2VSHy5t9KSE9s18zofwoe62lXZIzeeak4+cgUOS4ub4+MbN+yeGgqP2u4/Af/
0K102Ffff4YB7MZJVlqCFaxbWp75azSa1d2aH1KMHv48PXWTtWs+PINYIVX5yiySEDZjtCEOTWsd
H2W2LddnUO+kmS1CFfB7eunDZ4SxMO9F50qloWvljyrBYZs6gMapnQt2wxL2+ZZYDdDIeAJvQTNc
NzLswThK5h+nXHpraNeZY3840Uf8TDtM+5lB8RlX36AyEDOMCjPq+Rq69TWnNoVQtSpyEc5i+h+2
1Ew9vhzyqAVPktB4vGepQTueucujMDgoMTuGJjyKDWVrVtCGGpqei/dGGQPJFTTRhl++jaRMFnJo
0cqoE/tbFsn1miY4FntYY1LS6R+c+cbVic5dfRdgVJ2LBOUV1GyKS/MXyKcl9uxlKE5BXE5ovrA3
7HGz3qf8+yU3qKvTzLBd39IQ37aLRLxQL13ZeKbk0hHdvTou0aALAnKsaMv56Me1xFpiq4fZmCfY
U0z9674wZTZgj7BNbHY6EsQv/AAL+7qBznyCCWDBjyT+DyR50j44vJSeOWNqDRdnZz5qmM9oXqy8
tiktrVs/XRVcKp1FLTwF0FbjA6/fk6FLxIkObnVgskJIkxsdAYsnJPXydJbyFOiFu/wQblabTwMl
yInWiNPu9xce5i/cQEFHZKM95sI9vSG2PqdVTz9UGOBkY1POyQhZ2M58ZvyfYfIR1XCaXOnbWYnV
/ek0xVSCrrbYBlotBAt0rlovQPAfNN5gookg/+hzSepCH5CBZBVITD88/+GF3djp3Y9nRZEReSix
PS7oJ2KCTGOzGfyCgnUtxNNOk/Wfne1o0CiPqi/ydQNbo2qfcTf6IwMGvjxq072TMLnx6kREuytc
BZklmXr3v0I+62cMIn2GJrJK+hJ34w7wwGTE57GJ+7TNkNxVZNvr+QgVu2fHYrQNY9n5wAGky/Qf
yc08quXhV5hW6UUGtg2fCwfWvHVMR6bskKsXuv5/LWcwmLhpLj8smIOmry2z3JSokS/PxSVPeIw3
PuyVi5r34+lB4M2PXyXcOc/NZ0cM2Q4njj6XhcloL3OMI33IBSIeMvE6Ft1nqy1BTM/nPO7zB6Pj
Pw9g0M+fAOdrQRTCxPoHUA370yrsGDCwBj8VppTARdmu0+tmztaBqWsBAhaxBETwljO/cGUpQ56N
pN68rKcF27cwo7l3kOzh1UyAsppS75qY91AARcXj59uEQzs9QzNVQm8vj21oKqYkMgv9DPodV6AG
MB9DhZHSIT4TXYZhc2bBtGC21z98rVlGvi/9Z9VgamkeLLfykBvmkmChdsh4btvgXfae8imF5ypf
Kq8h0cK3AVzCS+uoBIGzbZ435Z7vsXpLp01iZF+CU84nuQg1hkstd4zgqfAoiVW8dqPheZ+h9YP8
3UsAH22Wblk7HWIGa+UORY2CMgjQrYzuadjBIDtvz0EEBXMLb2Mxvg3r5p0BUoGmefW9GvzXqjUg
MX4lhF+4sod4eQfPVoaq/h/u4DR9pVMAe1x/yyMRCMMlZm+63VclT+Hk5og7p9QTABQhmmXKPRPJ
tjGz3bRwB12s6htLJP+raW/MokZP+MYbRl0WFgk8e/Y9Uc35FWQLF1TR+nxnfswzZGl9DhtnT4oR
+2HMZzvHDsrUM+Q9WvgcHKDYcJLqZjuqrhGHU18eh+S5WOVczA7ZJvpFkW8xNLbQO+6fs+Te3271
Q51xFg8QubUg25NHSZlIYbIQQPq0iaCXZ7u+xmLCGP48YOrI7y7ob1tDFQ1tTKfmgwYEvX8EkrU6
nOGRtl2DagXqG2G5F5ast0PpGR2bTB+NhNFiVVPNpFVKVHlmCdibUEQRXAmFk2KC9CFDjicNWLQG
RCBOy6zVQLWD/BYNGmXzByC0CKmP0CaRUz5yzK2LxcxBtfhuCwm5X8VwRN40Jjq/E7Klonhwkplb
ZCf7ivIHxSg+SwNpKcFlz/Sa+FjrgPDUYogrr+KBd8p1z4O7dK0Mgx/vSDwcLocKjSWoK1zcrQ9l
h1QFYAg8TC2p0ZeDmVnTLC8HKo26DEp3kuLTMjwJMa7qscvBiq1mPc6iP/Ty++TzScAO/gcDXDlK
vSfhsR7Lw7PkCODihWWMS9luiwKkXliaSxl9KCKkwpploomOy2wjnY7BJvol7oexgw+hly9h1RmI
HbGt/3LdPAFjqjYhGyNTtoMN6GPp8S7lKSk4FbwtNP9fppyQLznCAb+h43pUB2DuHyuFUW31S+ss
hlYKaCxVV/HFepPTiI9SEtDKt3JWwammtsdZwFt7eEaC/cKerDPT2yA5jLSDHMhHmoFJy/aqYmUc
GNUWTeM++ioZCW2THxQ9syybbD7TRMTjHaIvWOJ+l0AUjvths7v0YF5SN1GVpyn/d3Ge1D1Upqok
b7apK9eVhGt8s7I4YEjCXc3YIyeXL6eKTOUnSFJANwatSARFomehdqC9pItGHCtrtHKeNOvqH1qL
dfv0Ni6KZ6IWa/zDhEVV1kkjHUxAkwt7pySjETUdUduup7XdroG0PXMAStsGXdzJMfdulMakuYJ6
BX3FFLCQm4HeSKYmZdjL+VzMT3M4BnnicmRcV+okwPFvuRV9oeRZvEEL+rtgkHcC0MjI0N83wzYs
E/4/DRU2cHytfX4/McLQiA8VaIf3aaY/XVO/jFBb6BkvirlV1TZqq7zKM/sTdwambYTV4Dndt4cw
oXcNs3JKAvhpeDN5sQtdT1opEO4usBrCnGk11KOA/TLSnS/VMO8QOEELS/1KSQGBjZ5yFwZIys/Z
D5WUil5EtcR4hFwKGLr+qswWOj8JgIu0CZgAjxsnK8dTwyh9INX7iUMdPLmtq0VA1RH6ps2D6PTX
zKt3Q0OqgOFHPUg/RRr3E0bNkPYNcAb5/p2rc/6ECNX/0JIfqzHd3ZFN2mYhRENraNp0PwuuO3eC
icAKFNIJJPXIAj5zXFgoGL/FVmynt/huV98ts/aBkLpU/tU8vEDa2sJYF9TMGVHRFu4I4ViX6hf3
2KCw29bBvs6LbIOOHXu8e9QnuSd3/6J/RRvtiWbuibKhoB+9DfBqKQXmQaxtQemXa8N9V2168buu
7d8ntcTJdRMjn9p78Y5dpssxOEhVj9vz9Z7M4yB5DGrKw1OhZQfipJE7t4tlL5tfoaMnTCDd9d96
16z7JMjJiNrUDhJiS6OeQfr8b5EqdnygFOh2Lbs7Rek9iUcJRH4ELP5R+a6pACTBz39bdg8sLCIt
l/3jJH5h9dlLL+U0c000CDgNgyimYKYsSMn2Q4PJ9a4MtpFIc9DN3gfF0lBS/LGD1MbD7sYTmoei
m7AYwdWp/13k2xXRUy4cEC8MDafdBXdig5zEcsAoQf/+mT5qOC1cn1cmSp3Sv+dlKLtN5sLhilLM
OqDWVtxhZnqLhLBI5kzXgARf3gZ73N9PDZTvUSrE+cdG6Pt6FYZqXSk5xRrnariDt1RUlhXTpmS+
eSLYuQi0K0+rM7PhPgHAYVtzvzP61sKxh8eQOUVtjGOzp4Rtg3+fdcWcuRKkn0qZw/OQGzuhzW8H
Jta3Fl5mBRNXCLJBGKCmEKLNJwXacwgZOmgmCRaDhGUdgC/vD9AtDCWLSqvEH4i1BHBytGaek7wM
muvT8J2q5Wu1TcGaJRoAlFOvvlU87ZhqWRVpXngxU+e7cNEy2iwvsQzC7QsLBQGdj4fZeOs7g7DD
ggGxKB3Dlp5IAKTNSE9LUm8j/45uFImXt4iEa5qVWF6o4ZRX2xbvYBo6t9/v2/kTiKy6o/OB6oIv
x3kP3s5zIVMp8U/8axnFsFsIDc/c9dKJIBBrO5/jSC7IWvvhxeHotbqPCt7f/rEj3mSGTIU3ClkY
55YfwyLd59We58muO6lrr1/zNdoEwhUXexQpaeLoUfZk3A6XdAOiizCVdbc/Sxrx/oOtGmri8REI
aNx8VdhrPjTLbW/j07cjwoEMjMsjArkeUoWd4Lr3wUHopbn3XjzMBZfQ0fAfcPUwgsHg7PZyNPMx
hcMk1/xId0/4yjrcYo9FUsxEeCiNPXUIik/35fJrQYFcoBCGD4uTWjvG7pHQuo/SYgQxa4MwJGEU
BMR/RwZL2hnQGw7hbpWlz/xzWOFlsYHOEzJygi5zDHbyM1/jZpW9LCMkDvCc6oseKcsL3GHZvTvU
Myl0++dG2Q4PuLQw7QWaFtXHoQWkg4t5KOTiTX2s7UqXS6zxuA2POX+d1i0sJYREeoYT7BXMsPtX
4mLWciunRhRL3YaFaRcYhDahfbjVghOQBKoTPSblwRJqpMMA1gm6afUJoPF5rbCLnlnT4sdEDBEj
BhZZ1LL/6IAPFtAsiHzztGS9doB9aP4QbqSmTC7BNxha8ifc2klztI4cMEDuf1Lenk3Wv4leD2ki
ldBV9L/h8HnvD1WQjZEY5K9fRbSjrmAcjVPlpPwG8SyxFXqeReOReq/qgQkE0IfjojaOyWe+r5/Y
9t6qa2aiyUatDluYVLFo3ENWvwfVYYqwF+rPnFpDMxcwD9SMSLqrf6nRsixscTS4dxNtP/GK7NcE
BIknGDwAx9nJoJNdmKwtRG91F9A70eTEqDpR97aaCj2OniXtwbI2MXOHTVyEoiZZQKIULOx9JF4K
wekczRN15jMoPhnJT7K0f/rJWAzQZ/pVepE9syFeNt6JmBRF/FcdRFQAZvjR+Xm6qPd1eMGbtBE7
1NI9mj3qeS5dBNn8w1vdiWBmPdGQ6xSVdhZY5xCTV7TxLH+ITikOcmZqUwjVBXyey9ZFJtFNBoFJ
RMwCGR+9kv/kfv6MicKb+RkhRbKG6pzpLS8hPeMxbeGxPr9qHR0hwhyufCPsjqonuCkd74zRMa9N
OVz+tw/0kX7ZXqiO0gm3f8KoaZEa+bLSQKp/z2euKOd9DmH9UJhYMgyPPuL3vUfjV9dj+mUmLFhY
gk3Dxwm0wbKz65qNcl5P0UjzeVQk+s0rG/TkopAHvJkEXwpx6HM9CRQ1mOq8by+AkD3E6E8oAqfw
qXZa1GDaJ9TwXLPUwOoOupd0Crx/BUXv0avGu0fKeha6arqUzuKOdl418GkuFVugUoHZUuh6E2jy
an8mTPvBOSq1FgQtWi/aP+jdgh3XxHL0wDcrLDjcpBniNl2w1JGn8vP15Gug2SiIoP2RYO8dQ6D/
09JP148FdU5QyAmT9c/VZ2ZapxKlbVrWtAiZ0rYWd7MuhM169vW/rVUfBLgvJTKGaoMj+CbFKFeL
oVbiz0NqDtziICcjuPkbC2Ozy4R5MsHQ9N3uIImXyPtvViEIKqFa3x4g3T0lBnWkYHPZZDVqJjaY
6ikRKCmcPkiqlBBXwH+2d5dBcxN4OXVlU1GouXNyDCQQkche4ZPnyhAXEsVlSyAH8i3tO6O9S1a0
rizpuUYjUqO0hLI0BigwceOhSftLW6ZgC5MJfPV7JI0D7aQ64hOEuV8kG6ZzvmlX9RW/0Rg2H5M7
MjP1YLYijHDsdeBngJ+KtvV4NQSGiQ3LKfnpvvdEs6d3/DwSa5FX0OuZZRrYt8FsweabcODI9MMC
x7Xs96DEzR0jxKOa9qdhQKeoa67nHafnjsxGP2XSKZgZAml9RKUJbQ6atDEtlN9k45oFdry9VphX
dWHGUqTOBmZevtuUjD+CP2H/ODklJcFjOCAIfWRdlAkd23wRwgcGwB7mDo74AjQ+yQlvQOZVERxw
YG8FIyOCfy6JtqpCDvzsHdEN3le5jV/Tmn2JlXnIcw7JFyHyI0i7e3b7gSUiCeUk3llo4y7jWihf
bC1wnuNAcZNIh1zXu8Dat5MMPArit/akx1XAHL7XXQhxBTH0BqEN6OOw8YGa/QhahLcZGjPVXMXK
Bc8SDKc0isrDLsJHBSIJYKELoV9ildBuU8AyTeg6kDMwST8y8Nud6VnMOneZ1J5H138kzPPs2O3M
cYcuNi+sFH4c3oHz+oAEjHEc2P/hPfFRLhVzdfB1qP30XplEvOnDGQZebSvrjxxhFdO0Ch0TQ3WX
DtL3Bnko+zw6kT0xMslomHyAaCWvOMxq4ulPbrf6/TuSgVH8f4wv6/HPNiea8Iymzel27vJAE6dX
WC2/GJEFzfwVBttwVEzibCx3wRQNe8EHSZ98eGtwPJOAuishhaFXHf0SZSabczn2zE4WhL2VvNIY
Q5/7Nx8+qGc+/hZ3FuFtyILZUNlUGzwL1JgXJ6lQSAPFWyLXw7CFHZRkYLLJ3092v79VnEbzyJ+E
2URmDPwFkWEjkvwn+1vgsPNhFIq0OqFjmwKm+Uo7VLcJCj0FsrTq7RsTGhKPqMhp7hXY95/e/cQq
8Em2S6skf/mINkiIFNHlLV2XfCPpp3TVkgL+y+eZtPR7K8eHPgVObPLYAghAdgegdbzD7LW/QWEF
+VuxDFUZPOUpS+zhV2jMFk8s7KHnV/0nrX5A2k3nCcywJew52ew5wc5d6R1xAGSwtrljIn9/vPTT
ty7b/VP1vyB4YR8jQcvp3CvM0n/MfNtB8bNiSwr+4hXdpwWTJmDyxvTrF6pv13YmHHEO+OCVKBmS
7VYvAEUPQx23HKZ8FbWNkWCFvd9HocN1K+kNXFASej8ZtVqbTvUCPpxSDVh1NkD6JgrS46856IBy
SlM/3kWsguje8zGqa5Afy46tzGmfk3i6kdOgAs+p7CZEGc/bJzmM8F4awWi8eDnSnAmAzUACqmf4
+Jpo5CS9Tjk44o1RdxPfCQnpMQcXc3tAymbf0X9WH3FCVqD3gJlGVHeqUgHZH400gkFWX1g90pza
857Lt0nREVVVLEjnf2j9PB0J2ajuH9l8oWbJh5w4CvniV/lPG8xRv1pWoZgA6pngfcnjdhMu51Bp
VEW25vz4R5vCbt18B8+a9rarxUJImZ4KEBHf9iLl19R+Pjc9ivDgtcJ09eT7OPYebcFvtj9ShrjK
DMI0TUJePugnunl5PySWJPbPib6xuU4Q4TgxFDR7OrwOBeQDwQygko1DZG/Ll5dcfgqz+g5Res68
/LTgJ7o+SgplQVZSCjWlHNica5OrQtq1t1xq1nCKQJFC3xR5pF4Vj3T8TJNBVxIbGWslnVV44Z4E
Ao1c5ul2QwgjpB4HdErwXnaWJQ+zfovBiG6+aZHW7iAqs3u3lb/QNIIHf9xQc0XmnMx1GyUYsKC9
SJsEFLDFjoxzASAdHrVM9brPcKWmQDbAYCfqJoEpBGlnhb1EPy/4FaFxgZGq7vywGVH0iydrc3xh
CZw8fYmFJbKzHj0CcuKNJdJt4zf3j9mpGQ0tuCNnAwud+ju8nu5AZ/Hm1X87c/+bDOZHMBTha85d
oWMwmJHxxhbMjMaeal/j29J1IRZiedOBQfRyZrRe5b+XA3+RgutU4FkNizq21AQd+WsYzKaOPG/T
eLUKnDInC+a8INMAGPx1Llmuo2dizbxr5IOBS1M8kNCXjIW9yeB53hNR+9WwRo41TmyP7JhiXmHv
AqdAGN8tHJ3Lo4iqVPPqx10TiZ7l1K+NLE3vLyw1wnTt5op0wm2s8rnVgajgswQ6Dx5UgTnBbanv
pF6eToXyff8IB2G5UIVn7aXyZVen6VL//WNAQCfK/tS1FevbCVoFdx20j7yFqf9bqwduquHpFHsf
X1SJUOReofMy3fZn6yxdHo9tE/Q+yq5fCwzPywi8IOmDktZmx60WHA0Xy1TjOB15jrU5JPk6E/pt
/NXWP8t950r54dGiDujV16kbEc5acgZxXbnBeD+r6dMR3/ZO4yGf+5Fn6Rs1qKgStUJsyCYB8nYR
adpq2FftFxdODAsBEfAyIsqxDN8Vu5gWuo4JTpJJ09g84lcvtqrnDlXSMbb2H4BCwaMY7digKyhO
9aa0GTj5SOadJkGSc8IZ9pXu/Bb8CqEmqOGHNhbQX/+h/xE8oAzjMnS9jCzocG2qw3rO9hEFNd+h
mfrYNLxj2bxhWFjgFv4265FugzAoj7YYW23nj1NuloHhyjQ1OKCrvlDxznMPfGUuyoUTE/GsZD1G
gxyUf5kZfwJKmZKsDEe/gKTv3oYQYZLhwTULEm/Ecw8Rt2RRWqIckM0wNrZOq4bnYhtP3kBLlvmX
emLq7Wp4b1IM9lZO74KBQvb5ik6FEqbHBVQ5vKdULf0/g0IqecHVzljq9vudlnO1d5ZCskjriZ89
0meRZHBkfcxcuY9vvJbc1gtL+R3ebu+8D/2lBoxRWDN/VP7L0oToV2RQzTvfrGsmH/3tc1RQdmMD
ChBKTZlDtKhPIyeOoO+gp3gP6PHv4th5cSEHQb4ggIhJugAixzumnGbLRJ0nJVYs+0I7GpslRH8L
ckqde62jyp9pAgm3Nb/GgKvQjdAiVmm1sN5eGP+W4IKMy0qHil7PIAleqdy6BX5SeN4QXsFacNpN
bcj1glF7ita5HDJoBfEZCq2paUp+plhCqhhXuI2VfIXV2ADr61oGOvBHx1GTwCiTx7WDb9EoRKeg
ZxwFwRsGSOMzQPyFBkdTyweRXw47bT9S8mxobxrae9rbJMyCn9SajOYn4QKumfKYVxcPoGa8g3af
CTDj3P1LA+nEXp7hUnZG2cWjTslrCPPBIrEM/NACTNRezDh57aOaa8ESyPrpaQEYm0HZzBYgxbiu
FLFcOcA2AOqi4x6R3190qbfG8KPjOyyxQEGG0W7jmpN7+RDzTdxx5aeeFDVWB/7xZXy7ifOiXUUv
WrZilDGnSrz8wBmj6pOCC7WJG3/Ng7QzwJhd4GpraCi5OPpxEbAsXnuoXf7uYXVdTPyTvwxOiVea
xiduJuV3bDAA49y8YB4t9wTxg1zkJrYD4ooIj0WdiqJMvGX2nLctIa2b9SpoWIkmfa4GR6T6i/Qs
15JhSjSv1TUSJiZnSFKx2lWVs9APBNPen6qNE9oZ5SWZwb/XnSC4+JRAzTn/NpboYYCJ8PZRXGO5
jtX8V5tWwudma9UP1spz+dHkq4Zp/F04n82F+45ScvsDQTvjCHKicp/qpx/asG+Yc1w2BXxq635K
4Jx9JAIJ4YYJn+u1wBIFQ58yG5YoIfHSDs/ymx8rRDNhrnT5/Pt61V2Wktl5RV0Xg2eUziOUkMGI
qB3qDt+BcaRZtw3vZqZZMOW9r/1Tb6vyeW+gD2d7FaCG/DUYB2bdlr9GHvdLFbc7ISk8ICGo2hdu
fyG8SP9x4UPOc7fgh3tAFZojDtDQ7wKpykWtN/2c+zQfx9pS+sZGiSb4G1jA4kBtYzmAoC28JU5P
03yXbJ6k0EoGScJNI887ebSAY1MwhcUStzuhDfmyZ2Y8YBsfDXErTeoxnZP6CqERC5st4P/lzOf9
B1omX6Kl2QnumLbjKlM1ePMdfHui5DEnxgLoR1OtHxaT+ZfdGc+1zlHrJJzBPyuRAGO2qx1FAS2F
22CRH6sXhLH3Bh9rudh7eWYKcmW0KheiUVGnDYUTupnYXOdGNPU8HeGcTzuqpn/HtXKF0EC70As1
3MfZ8zcAohntB73dfPMdyEGUttXUOapPGZZq0W1S5jQGnntZHr0FJkQNcJzGGOhyzpMDovsK9bvq
aARa5h2EY6opnXIGDYQUcheVqhYN6L/BW+Hxy1D+lKpWiQAa0QPXuXLNK66CMe2iH+I6kLiydy1C
6AXil2bUJcHwbq5pRHK/O3XpBzIRyNt8z60Uv1CgRvBDcl1d1Ko47WxbY6mQV5GWuGvyR2RI+R3M
XVP4yRRhJXoN4OuBMvhFjBPnOdZG5BZA4ltEtmkJV37sYU6UGV4NdOSq4vyE519pB2aoi9omftfW
+G7bnsWVScEyah8J+YvWSWGpHxZ1dfp1f5CI6KqlolkVfbb8aHaxuT/F0DD+OWQq7zVFl9dHBmi2
5MArnLjcCZGfkkgh1hFjHLmPBQ/+ZJVE8/hKyTszsnbzfBv9o760D51g+oLwBYrjFJEpgPXXHOfe
tEUOK3ur2tcF4/kO1kc07n+nZLEXroMlyRCo0I4OCUDfa/ITEVpnzx/9jelY1LjlARlGBrPRPJvC
Txabjp+Evv9/apqr1hmHuC4NJ5p00NZkLRuyWclKJmD/VUUnOkX8RVQR8WVsgkTmuexw92St/MUG
KNOh8hXL62rsIHaS4hXRhTOtyHbpEmU8nhEP0GaDq3vhw3hH5dwPzM2xhTTSbTj2aaXWaAhe/R+/
ciKJ0ArOhaLpTTtlmBv3BfdRiTP+FNpCsn0PAbYRumt+0kOht2gPX7drdeoQNW7M1zzTOIoulnL1
bIWPUZKVWxa/GPVNCCZKTrF8Lmtm9FvXJmxE10fE947Ep+/sFjSqV5iRjAN/N2rEEDsFEy5F9Nlc
Tv/rJsNYRtIOYe9w4xCRL7EWIWhBDDOWsbQQJbCiizrZuK8VX06AurEGqHy5F1Z0MTZ0Y6cdfoS3
5Pov17G6TZ0tHFLkx2A5KGr9ufIhabtBEmDTuIa3W6jQqt+EhlQeiy02FEEgMgRq/Js+LWlsJnhN
mYLkIKOSrxCq2OyL2phMFNlwI/DdCgLTIcbe3cKbUmLNt5Ch5DPvK4QK1kW8Tmvtj/LP+D7//DhJ
ZRM+WzsAGBSN75O1nko39tGk32DLb7JmYkMq/QTvtB+vgWU6nzecO0PfyiyOy4VMiw+RRUIXOepp
40SA2TP4hLWXxGxPKc0q/wubqYCwjJSpqGpQeR4T94pNrGuWItu7zvho6KhftgGmPjfAEshOpjaW
zinsBecrzPJXfj5KA4dbBR2ZVhuXwNgEx2kvcFgVHOgAgOH4CEIw1jMTTQhP/MuRJKbkk2NEIcqO
KdNAFdVSCAQ6f9jKwnagvBcZVU8ZKAzz0RJ37Ntm4BA2u+EVj1ADKb9+bxy0SugaMdetLZYAbvBO
7QApGXkO71rZKu4IEc51oUelTl7QEsUzkjI8GheooYZUmPdUlIB9bBR5LTmYPP1Se18li0mt3T/p
NqFSfs6qeFnou0VoD3U1pPfMbsBCqsJocx7m3IiY60I/wjaKSGNDUU3ihPfZejL8LxfsIC8qRiMc
MivKxcKIBYprErvXKc+s/AAtK4KhWQFsuvdCRtFPGgKoD/Xv2dsCJ81FbnbaiaifkAGDKXYQN3hD
EwS3CeExOYDIFKwdB/TedopMhYfrUDF98J6G/evH2yR2zXKReXqxzH8YHHywVlAW65Fme5Q3jfdp
oTOXavgwXNNEhrBGbIxH5Et9BpQkzPBS+BYg3w4zy54uL6tlz0ovvb5av6YjDTJO5D2rqUMZ3A+l
OYX7CJXvGwzCXI/4SjpdNS6N9rdhkW6sWxYFPjE1wemlO9FNdY3zulNtr0mawzB0GAIYZXg7RB1r
yPSSkSu/x8SlDZbeziep3XoZG+VozpXwx13/qDjWezjd5skDvGiuIK3roD7a+6tt949YeuEpOrqq
9Ftngup+3Up7bKjF4Vt935IAS40H+fxdyqklPUkDwggyrd/pLnMwxB2CMSak7/txlrOi3WZcHE93
s2amq2VVDLrSFW3Wgo5VQuMwRsBz8gwBLg5F1uwHD/D19gSU49MLo9jcd/2yI9qpNpCBI/H8QAV+
TTfW86PEfvnIHxlyEbf7s/AeAx/TxfPYDVnXHBr27fOf3yW1as//ObBY5hRzGVsESlsKEunXot19
TaaD77nAx/uoTOeIaT+CRjH1tsAe+FE5U4swhV3XBdcx3IIkdk1wdi/psKMLE7X6CH4lbX5bi3RT
3+1HCFU85EXUTZ2vMmADIR5fJOcMu54XQguDqae5EwbBusVEVMhqAZnK0M5WoE7qlLCATrQzvbDM
06f83fGPCx3q2CjJwOySrNAwk7y3SmZUVsBAGU+hVfw6FDnT6LQew5hPdXCa0hI9knUtxUM6QM1P
7+Q9x44417Y+oFOPxhur4cKUfUAaLeQ+Te/7d37F9+pOwpj0E2km3fsukG63ArCLHLToRaU605uC
/+czghgWdHBMWnx8FcacWalO6UCjJr2FWLMUHikEq+50R+zZhVBNAz2DtHMndQdwgdWDRMLhnHkH
Yhfog9meT+rFsM7VpsbumqSSI9f6PWzlun8owZhdVmjXe54rCx8AK5RGrh/TjyNg50E9WpMBBSQ5
eQExhMfnFXKCxdAY6VgIjbJ2aP8bfIHw8Xb3RNb4VBEdlIDTqndvrmeVVaPinRuO0D099GxS4fRP
nk9hb4UaF5TWKH7fWH07fJ1ci9snKB6tJN/OfMufDRoxtIfh1VSIHBZ/dNafvrIKShdRODeNByhV
nMRmS9zMgiZsWrT4A1ORdigO8HMSeg57bDGAM1+jKr8FYOmJFrgzVOM+EvzfT4h/bhBLTIrRIwUW
W8+ODPvvJu/jeHFq5rL1kXWZhf6LjwWeH/B+bzlXByDxV2EjE4iEinHuZDpDe0RTjXX4+74sLUrt
BYUs1ic4M0KlRvFFCXMJMZg6I3ThoD9XPSrBgTK5tVcD9d4Ql/PQFUo2Ip2tOB+6bsuMwlmaz6LF
1vMN3OW5IKoaQLsGoH+aeWT/ZQepPnVO02HgmxunWqlk5yne52Kb5Qx1xTzWqywVc8DfqdYN1XmN
08u/C2R7TceFRrRO/FrW2fZ0ilbbLnR5B3sP3o4hteCEdHio2aSD2C1foLc2b4xFwq3aGIbomIZl
AgNM1t/UwTZq9tGUB2NWS/HCEbxRXbXArwN+MGcP0nJU2IYV+nbF33NuOADosMG/jh0pF9JtEE+X
Gz5JDTQpcC/iHCnU7QzowhDRYh0xZnZGwqjfKSj11OYCWa+oNG3uBjn4O/cqTT//xpKZmot/noWc
g8n9XCqaksz1m6sGqHuPgc2YM3Xw7vHT3jDtxZsezwj8Z6/ziyw6JDsENOFgZjnLC0wnZjjWRrmZ
vgdy0V3m9zOJtxkh1X75WOWxVdrxNrzxoSuT9kHSRR8jemBDxlIsYLEO8R/BqAtJbHKtP8Czn1aD
gtX3pFBRtyeHnOFC52TTbcVPzfgAEJDpGd/4faFYHpivoFDpo9Uoqr/62cHeBe227VTUWCnhfWW2
ApepqsXoJQHdD8ar0aPPuuSBdxMNCEG2o01DViSTdze0IfPC9n/6YXaMOID1pXnfT3zI4Vt964qv
dbs5NGlxUDzrxpSBVhF74uwJ7moo3AcyTHEuaHwfMA6rHR93r6hEaopumIzf1mPZACSANUMck/I1
/NWfNcfsciGYhdubCivtrxnVUeOqrWu36ZsF+1QrSQ70OUoWyjkFR1PLfiTDqFL6PrJbb0zVZ3n8
kNDk4dGrvSsSW+NEl5/LgcxKRSIqRXhC4SyjPvGcuJaQCOY4gcOpHVDKwlDnw+kzF9ABT8+DtQjY
8YEFHvUckcHvvEJMV8rUkcEEPHZsRiXupgibWUpKhgHGq+f6VQMKw4gGDFaUlnGblkqXyWLqiGrm
MCgPXIhpK+Z7q3QC3sUhh61Le8bGcEjUrRVKD8WAV+OsmxfQvD/cpPMStZ5NLgSIBqNAM/5x5mo6
IGw16XswsWN5EneLcKPNsUVY2stAo6TvQEdDeLDm1TPgFgZEKsQnEMcDkKnnvFnsacthN0rsmkHs
jE4GFOAWLoDn04BRkO31/teTJXuKa4FflaaCKv54kxNAZsx2c2kiMkIIoZnjQgUYdg+0nivhMrBx
WxW4jvKBg0stpyCrnrF/7ZeOuZ37wITwf1x4NM8HAS5o/YLtYkmdb0E8opb0KMDUD/41uu9GfUD0
TArrf2EIsbGGLS5VEsnegLWS1ZMYEDdqRxcEHhc/U5SOMn5ohJ0E/xt48b6K8db6fQWx9q2QNM0A
vRlZd5EDYE7vYqJ4Y/SabUi8yMPp5MRqTTmTnt2XICkGHz4r9IkxRKug8R8dSn4bQJJrMlQlgx+E
JDJAb1cCayz5vQcyvVa3TVVhw2ab9LvXHusXZWHKJ86exybyqesO+0+pAid+wJWtjXM8HVo1UZ6/
H5r7Kb9CHJ+3WzEXpRf2BNwL+LjuyxrbM6jnC/HWGUk1ZsB4QRqIdGMj1aYc79ffzJvWtqJdKYda
wqFyLlgEdX9vrjQmgz6vrXUKF07guNWkZf3OVG9v4BOAhrsFldiw0vuM0EjKoJg0XDLz/BGXR0Jw
KYIWyfN/d/0IFyj/XVAQ6CcTIPMrq35bOHwbhij/xe+uSIP2q5OjWbawx1Oi6N5piaYhp7OicHCD
+E/pxjIz7eATfVcI2P3+LmoK4mZu8wzom0QRdWLKj+2J1+YqBS9BbO8ov8dSBE1XFSQIZGlNFuRz
fXK3bnLofcGfTwkNbTvFuvkWjymDzdABR0Fue84Jm0BTP2TOZF5CURHS5MNntQjjs44rq1nyf4PQ
+boYGJoT6k6BCal+7WWPp7UNXFkDK+tF9abqa1NCu/vf8qbJqaOMRVO7Sf2W15qinArJWjISomLH
mG3PSR3IAjcX+2vF+2Zh815qvw7ko+sVYYh0G7gjdYfox2Bd5Xrt13G9IGnpIxuhmc2ElNg3aA/C
qgTJbTQVtuf6MJ0+s0TEfJI7UwiWD0E/RIFsF3h3wVXsZN96bzCWV6w6Qe70bOaNL4UelN6bvKY9
VM+izk7dM8NG89nkPeot8gYNnmclOHUR0u2Mv7AdmI5f82n5yNrs/Hk1FGbe6ctXnlYrP/2Fjl4j
mS6TG85XtWW1qzh7fOoa0fg6Q59berRXW9lcvN+TiiEIpCMVhbqeAjJeQh+zcPIT+Yfsh04h9y13
98cDblxAChi09RFipcUCNvbXiVAjbroHx+XPxV505AFKEBs4D+M2zw/kXvCtPNBWmu+WPYLvJZw1
tLpZqhA8R7m2KHBni6GSJ1pRLY1Qk/lEnkk9iQww6FQacTYYUkMG16FuWBM0vPyavZT9oG3bFPgD
I7rOTp8LSTuJ7TFVt2H1+zZ4/dqYnetAgQZRmnJ1YMqcIIyP4V6ibzapBm5Ccwx8VA6+hdT2lsJe
uWUmx4/fdVbTnpz0N4zzC0vyyd6gGyWzYniBkPEx+Pe21mcLE2aX5jpaaZP2udlo98e258WX2IKw
5otHpXCKMarJQOh6YTExTTT8jIXCFdM1rqBCtzbMgkXM0lYspYyLT0KFREZe11ShlWMMamjdChrY
tm7Q+i6Er4Ynt/5QLNjhH8ZSs4BFmdEHhVZw12LeFDAYZjonAlCSeV0D27RnzbNrDWfJL6hSTeqo
TnsOcu/RQaHN2N73zFDr3ZyZAB8l/r9pas4j2ekQJ+MjAUfyuyafCKTbfWaTdoh2Y5j+Tf6lsHO9
Azi36WCQVqtpPZKFO+EcApxLVA0gJMqwO2Lm6L9x1vIgbq2b23NfjvmMa0SAq5aqRUvw+NCaLg9q
3ClDBLRpkFEy+E8uByMSLo1dFXy/5FB86i1c4gLdjmhuMJrB6sk4+0c/BkVspo3kXseVZeBeK3UV
eZCOyNgPK+cQkVL2gbU6wZWdAjKW8gztvSM5+xOyXSi/MxFlUqWMAYE9QtPETYGdGeQD3CU4r1kR
EJZGa+ZRQWJD1bi1ucfON4toZEyPU+C7gGmaeBBKHDzt5ZDkbE8ihdny43OkgssPlv0gdrhwE6X9
oPO8dUg4MlR7zkJzqc4Oz3HZ4dRrzRffKVrW/n8kHJ9Vn7NHJRH2e527J2z66ymE9jiT8GLv0OTj
SHgldQs+zYrQogXPqqsnZlWsMDMMT8geTjUFneqOqO07LOKFkkJR27UynlPQw4pCZt5+RsFubHbJ
cu2QaVJu7CHrNPk5leaMC+y8aqCmgFKywGe4ORTU8P1bJwU35OPxTqk2j+5g8CO+WUTXjTuMiKa0
ZIZPudTSehNFthUbHAOv+CTp1PRIaDS4CvzoVg+oP2uXol/yho6g+pgyZ6pGQsGar3j5/UhXDR8P
12iBfXRNP/PdhWUALQuIeh7YB0roADar6Xp33HDLDCBkv+AtZnPwvt4eqlVS2tiviAfIVDviFQ2A
XKdh8IclzHel8r3neXdJ+9trhyTpg+fQi4/o0Zf2c+bbh6OBNhLu5Y53PS0EidIJsujwmlO/I5lZ
mlanIvDrprqSbWvtQ4/DFP540vgdacnev8XewYVc+E+lqzovAemvbre4Q217nifwaBbwds4tZaI5
nmdJfBwxP6PBmFFi3dL3g6vvTkbECkw/hAM9CVhHmPQi2PWIMF69sdPoGWuNW0yiXZ9OHmgH0Xts
ieqFhmf9/m0ZaOfB/1BpC+9BTdlQ9jbaSbINWzmOy+vhfGKMzOCJh0mLl7x8SZPCMJx/Q6KKGrU8
RC2/Plj86Iw1V/kcvlx8/HGtJIPtg1TkfEX2YywkzJ34jw4VzRZgPjHG6ZJGtYoaw+w3fbill0rV
McdKEWS3PEP+aQoNx2K2WBh8enV+8DwpERwoNMcjHjnF4qdUTLM1VjQbAuljVaF6vlcSWGSbTfsG
w2G77bCSBmKQWw1TwiHeInWypAevdTwohNihBr5HXX89ko6MCt7GaAwJW11huX1jslT/P7m6t9Ye
X/IdWctQKUV+80rElPMjQP6mK5O2cnusC3+4ImbOKvfNGba3F6H7LSrJb+oXiKhdvCIxNycU2bKX
b8e9fxkynqp4Fuwt1mUxqdWxU+YeeVl64ZKuCJGzMPneh5v4jDHcUsdPPO8QJNAkXZyHoPU3YDQf
ZCSykzdnUiJ29pJRj+ritITdDNZCnPE93Blo5wTWg0+AWNi4AtQVMpiuqb2t2MNSNLvrXFW2IABW
CUHlA25sUdGmdYtILjDIHuN/Kg/5XHOI7HkBXi68ZIetyO0dDaBGLLMPrJH7brak681Qguow/axv
OuRjzyh5au5jegUZz9TIwDENBwNlRObTO1xaJQZZZxeKv6JllPk/h7Tq7kl48FYgSHxNX2PMI9wD
s3pqHKdJ5xFnta/jnOS8I3zB8GJMUx85YEPZ3y+MAQhm/kzad5Xgv0fi84cbr5nDKoCFP3uZKHEt
6qkOMXbPM2R0zqwdPjWl027xGJznaTwKoTD3AGJobfLt0bNlZmiMWXZX+h1VqL8Bp8Yert907Os3
27sMw+uDo+bNfCpsrCOqHBClQd5Ux6FPszdBhi5TtKM3/7ZcbE+BJB0KLeZrqdjzYINW542lyYMG
If4cytIVybZLJ4OYJ8D5lnB4UXDteivaxoMk2l/2bsSJprjiN79BmzQQrOi9Yiits8iXbey7cIi0
EMDZfP2OypHTahiNqCgVXP/C/Ukxae8n54v7/ccmCTvKu6fEDcPh4nB30TZLjG7xeRSaENSTxbXz
92vSyX7qyir9jiAZkL931HTmwomJua45y8J1JqX9N8OYWBRw0sJ00mRyinZdJvkI/Hk8iGuI9vVh
fZlxKukDcfsFpsQVoBen2R9hv4XHg9+b57rBs6eT3FlCquknj5Vi1oi137lu9g4FYWNeuXilGO6M
veSw8OQCi2XXUoymJqbccVEsGHy6I+7wo06XV0rupYCFbNDtVyCZWmSCpjNv6USxVIgl1gJj0Qo1
YX0Y+MFBFLsA+0c7lhTGtLCLGgll09HAeD77THh3M4zLJ3tUgKW4Mte+BEjFQVXdhxLi9nLScllZ
L/YKISXPsZsrkuqo9xEATKrzadcv0Hj8QPcIAadE3HjcCjCbaGKY8WnGhyR0udyVfSi0RZyOmWCT
XHoUW/EfyL/opg/IUtH7LbC5y5giGULi8ED8ggGYgY/Soa3TDvVnjhAqY5k89z33J+668eWmEJdg
jgw2WBTGYI+WvO3XRSvmSw8kVeKWqm5G+k6vd9Yzjo30cu5A3VC4iF4UqmXl/gMJ/wLSioGfpQ41
3i/tf/bd1t2MrP6Nu5HgqO1hvPY/Et49LZ3mtyGntgxE6bcv27ea/eNuYPAG9mRbRqRF0AzznOBv
9yaYIJogbyTRdvoOg/Bf9ZuIXRfERZUjegmsj+/kVifZTNSgWvjLQ3Gyb3Pk/FxaHo6vZao+4Oh2
OwlS0p1mVjf6s73jvEKhrwYDmzPu0N1WvtE07emPKpMN9olQuCjo4PsHQkn27sS/sgbJ2m85Nmr9
bVGtL+K5vTp0Nc5DVXCcQ/SdDEU/m0V005GYaf2hsm883pjIiKhjnlB5124Ur4xBFuu9/LXOGjjD
VXbBeunlW+iAK00pxfPdrzsmitldAYGk/xW8P7fi5XCuUV7tcyg/dSsujfFiTee9Pz8ikzhYcxGc
leArEMr1ZnvjjN5STA1ufaxnmX0MpgDctn0fVvIcxossN7tBXZ3tfuj9NBzhSo8ckPFuD/19bgCj
L0TtpW3D25GcZ3SVkQLmV3Zw/qBltpr2FoMUASafp9J8We06y8Knt7iML+sU7UzlmP5u1JHrGgBZ
oN+Ab+T8KXkX3DcDzpkibs6PRg6hgT+PtS8ECWOGoQLmm6W4VeW0BNaInV49R2Q3XXLC2Na8Nqhj
ZZi+YjuFs9GpUwJhBCUgC5QNPMaWRlvpSjeiH61jvBTeLAB9rVZSNRuy3bhgNfq/sWFfUsZm7wJJ
ZYiwudvtFfkbzqcPYCiZo7EhJqtZ3ujCTSAZPSE4bivJM21+L+4q5m78jHf2+zkQqswRLEgdGRsE
UWL3yMSZDOCKqsE3ZIrNSqmiO5usleLJaiaW53bW+HZIMIcSCZWcNgDFBFayfTxKw/efDaJUEVyx
k/z3UZL0k/ONzlIeRMLrbztnooeHHYf0cReDcTSGXXVmDgsD7OJQTKt+AKT/IX9elLsYsvq16pQI
SyORPcUfucvVFmGxvZ2LtdD+/aok/7rIBHz3dfsadlYMiiQcig4hQXZyVf0O3T88qtIXHuuXKpor
5axFWjY9t+Xm70vt5mYsB7kwIjRVaMyjSbLNULiW2qi6kdaJISgBAtHvbEFpKT91oV/FzFw2ksyd
Qln/4aGtBhSG44p5QNq2UbFGgJW6EQeFNoEyydAS5vzafI00sy4fKz+xbcp9ilgTK8oBBzcESeFs
gOtkTo/EgIQXaJKdJ0fxjzyZ5etqNU1OJuYY5vdfpIr6W7zvt713GWIG8EJLSzrd4BXpTbhIbE7b
Pu4phy2TPw6hgJr2kZzAAPN6YgNaqbhLF3tKCM6xzSFL/MhN+aYYwDfufrkD2mEjv3WX3RukPIea
98EvnZsccO1RAuqSWVWNY0Vqmolizfjfr+F81M7TsYHkgq7vCAxbnhzVadR+WjrK5jKd32VP8uEw
YF9wQOk5ohLGG+VNB3/738gS/mi56P/cf4zC+aCrTGPoDVaMf1K5ivyRU7NXx2lsoJTW3/JScARX
ftSeDAiT22zEjxXp1nEoF6XY2KNGfnclle1w7OjyocuLE5o2IreLzJa9Toh3ZtRt2ddomLIy9u7E
2dj1hYUmoT8jM2Um9OIYcnXfA4F00+ijpBYYC/NcMCbCXVUUNjDeTeJGBONGTRQfVDpM7dcF7k2b
g7WZHMVqljLxQFMJKTYTzURCjYSNN+mH4B1xLPA6/T8WN5yHjUa62c79MLHhBJSsSphturpw78Vj
54V+Agyxz/GzzszlYZvntGdopw61wB9OrYLeysAx+fd0DefoIcVYWiegG9ak24oFrd3unSMc2LJu
NSrip6S+XrRD2BYk2Lk55cTtnhmsWjdS3iVUnSguUrc2KmW16IMa5I/6zJYj3NSam9CcqFOLe3YT
1My3bPRrfkV3oSF9kSbdtgwPBycM7P+hS1E6+/TwZNHFuNY66IunZSvmi1Q7MfeUUmBzzzN0yAMq
lg7U4vfKc3jSMZlsqt4z43rHtmcq2f97vwBje5qSxkxMxTYCFpm1aDK180nMrF8c7zD447VLb3WR
t1rBOePp6Gs9DSzAd17/PRNIm3rnPdcJOFDk3g5P9vw28FmnN4Nwg7hulvvx8mEiImLb+t0JlkXZ
JSW+2fx7fTuXuJ1N6+5Q4CgdAkrCBMODUktoff51VRqOh2TZxjjFfJE+qalIkhoNIcK5AThuka7o
OXeJ9oIaZe4/59AIDuNnxii8BbXQKq9Xg1i9gi4wqDEWI5UGkpW76t3td0UVIpaTwpbeyjheibVA
7jmxLeHWpfJDvmp05L6FsfAFIGfGNhNYpY7pqQCqbDjCzV7CRh0avPZ4TlxzsZXBVb7fvnJONP3t
V7IVJev/NcFPT+0HmXhkEsCQAzZ4v66z9XFiI8H0mVjY46s8vFdlkC4enylKwSzHW2IcH5fW1ir1
qM86OLYHnkXiOYEH+TqezcX9ukXlJL3fpidy771RCE1o2NaUgRKPGH3NUxKH+ON/2PWecPE7X2/c
Bbc/Nl/2gm0IVlujh8mgLuWqSIZSOMV0eYHfPXDotW8WAGqOWPzkTkhTYuEMr2l8h1tN6frKsOVD
aLzk2dO0lQa/KDfxREXfpqRfuZJJpXsLCx2PWTn2UfAAVFWmRdLFDbxtPjB3n5QIxADb2KYwjuRa
GHhLfjIthKCLW2YjnetVoMCD0HvUeiuU7HaFf7pWzF1rTzji+fhV2Af27rjV59uWsZzq3geKjybA
oc14jUad7s8dzsnLlsK1MKU/fx+BZa0AfqOuSPigznQlQNkGMS6PyxwfrVA/3udTRugnDNoUsG+L
7fyYWBPPCJxy55hwVcQxwK9s4qX+4HXu8VGo9Q8J4ud5Gzdorp+JlrVfSUYs9rehgyESj8/sS2ZG
z+hVQ3xyNMWWGrnCCKMdwqT5aU23IMJUcNj2mdvHa3Pd/0kV8APQok+4okUtJfPW8p01Qi2Vtz8p
/AT0vVUu18tGunfn08HgLmatSXeIfxXsCa6w/PnWBaUY7RH52OldsR2hKEB++8gQaghIj47Lpkyz
v3Ta0bm0ZkvjG96y/yNwT7uwpiURF6bRUufGDqAtuNnF+35Dg7nsS+EEP48MiWAPJ8Ecl1tsV6JW
J/qv2xnOTZtU5LJaTqXS7dx8JfWwfaV9DH9mIiU9E6eakBmbNYFbgCf6OGEbdxA7GjR8ZuaWdebX
sGLdOk3XyY/fRg3lc+TxiHqDkbCDRtpP178BX08AsfzJse91DsMmd/aR71zKOqj7hamUbIcr3NfC
LjKW1QexUR+N/vpOqt+vXievMrFLOozOzoHPtH6T/sxMW3cwJiY9zg8AoQ3ZhoAUUUvb3pX24FHH
qQh+uJZ65ejH+DSKzu+0dG+TKFplFxiY7AXMPBoZ8SNx7kY0+rHfE/QxYPCh63ohhWZCALRuvAgC
PB9JadmhOPbKXsewo0HH+82MZi6xZI0MXJzvZnytxACdZ4Mp5gCvPS6hvJXA0D27dm3AHarX+Z/Y
0DItsPyATvzb0JeGIuCrIlReR2ZmN+ESrqAVrRytGkXQJ64bsEBQBhd/HKM757p2kkXL93SP8AyR
X37eLrxqSjWdNq1EMQ8unPYSYo0KR2xwk08MCRIpVgY3vSY8BdzokMgkEXEw35IDP26oZDa+KLyJ
9v7+7GvvCQD6Vpe6CDAqBokcV2B3IaNHrTY62ReOBvyyiRdMCmIOFQqtIsCmb3t+vzvpNbLe3JCE
7GNt/raDm34h2E0PmIB8nIiC7yaZ0ZisrJs/CfrbSJzm4YHSbMavuckGe3v6r1YhU9UfcgQ1kTHH
dKUcoanQY6xfVw6XLWBYl7g653hbxTUX7OpVjGn94r2iPzF024seSRWozOTCjdZvj7+qswmKOdb9
14dFGo9ArS6TV8bUP/bq/D3/2dTC2RTc1ptMYYe84VRBwchnVvRj8nO03Y8Eaa0CgvWg4EtVMMhy
4RST3xArEqvGd6vH+awphcY8UaznIpSx94WY5ZXM+DLoiX8NBYcK5Ie/72ta98LRWuzPB8aSKTdZ
ZkaPAaSifdNwQa1Vy0pTWrMSBgU4bzzXB0cAwZ8GeTQmpnua/x8GCfY4HLB3UoibW8053F7hLlxW
LTbtb5yJ8L4KqCLpxMTw/M6CIbtYBwcMWwi3KuXnMbYgd3f1y7VZu/xe7zK8UAw7+n8Scf5miK/V
t6jpX6sjThyK7zpmLBptb/XBe9KYQrirraf0cTp3vncnguVoRE1LOlOFh/Bk6icwTS3rDBQRBD1D
RvV5K2bXJ8RJIZNGBvtlD+OxQ7gDFzx56wJJJSvRTsa87J3VqNKzZEMWnxb4FnKBXc02ULYAC6Rg
QKrGLAF0GuNqN52+JHPVGm4/ZyZ42UYeuu4qXmO1ktxAesU094hdhd7hd16eof+2gY2E4nakrUn7
VrdGYjRNj6I8b85Qf4aoEuojheOXpEQut29QnM7fPun+CcY1j7zbTJUlhEQsw8OsrQlSP6W3td9J
VyJWMWJcpVxmUGR1X7C+TWDlckL8L8GvVtkdt03yLqkOVMQb4qWT0L/H4XXdbl4eWyiW3SPuMstk
J1vS4HDNuzDzuuEwPFl6oKXirJMrfBOEx8co4Dvu888L21HxG3hTF2tqQaw6vXXIAruUkSSJmAIi
R9V+vBvvuhmXfesmb+9dQRM819BlrAAm0V8pL36diGXc4LwZEevIsSopMBqyk+IqcR4RmApCzt4/
tvsTb55PO1/R0/u3hFy0Otd3Q+4p2vlX5O1PpvhYzc/6rH3f8AENi4LA7wL2/oSIiXX6gtrpyKBw
kOqrCatYc8y5K6NKs+9tffQe65CBWwpvG4XGjV9tjCUZ8GWUhDre+y1gF3BFJx5TXyo+vbkJvXNG
ZeHY4JNgkBuqJXI+xVsmz7LJpp9TYfG/3vBl3GLUuX7I9WPdX6U1maLAZHHLRm/vS+iEn2277WUR
ylTYoDDUHMLvQz4Vm8nzrHZUhFeuC7aF1xliyV5xdjpDBC3lZXIN0R6jq+1qVNiFAqFRSekDs0Yb
LycTjP5KR3xMYBlpMckmgmYYWq8YppdsqCd/9j3Q2R7wlwp/SM8GckRSdkifM/ps3rE8JEZdKQQU
Ft6c1Bzf3p7dtMIWcEpbYTiKLU6q3enDicZTt7lDQhHEec9kxJWqCca9HuVG7EFbsBVB+koBZzJP
b6mozZcgidNvSqLPvI6pceNcQ/EAinAVpN5nNNXxpCVY7qRsffdFnWm892SAefinStcrR77B6gGk
J+HTnnyRaJFnwEPKjcSHOilJwChDi5VfwvBEIoluWN3QAzOiBL2Wze8CZgDjkFOEzBSQDRd2LqEX
Q7EtQJa3BZOqvK0L46/MEe52ImjMARF+oMF/hzx9IUJsmXjcJW9dPeSGY+7pICGRBpHyCD7LtRTC
8us3Vcu58PwbUPBw0g5ghBZPzEQBuG814sV/XvXyUzSxLXQzTPrWT+ziDF6VRa42Tp/sdXOLP6A4
lXyVFh67PqqlyLFlEfKtzJek3PGX2xZ6nTlq7jxHbEJL/0mZq27T8RAwv0QLmHkoVKY9aPn6flOL
gPsypTw4yqhgdOgS91a5WKCuFUFl+NNt/h5WLgeaCeEBVYgnn0f1jyJFyrUy11s3kgGtKjR3x3dX
jJq7cDtiA+0SF1Xy0PG5V/G25OWvyXc7KCy2zjdp6Wctj9ae8azR/fX09MoFX3KKt48IJ33O6nsP
BhXsRqdhKEMlsq9ChLqIvKtqKRoiJIGkuBUtz158e3c6hEkFxw/F0CR05IQQswrfRTh8na2P9zWq
pgfm0mcg+R1l8aeQdQD76KKBs+ebYXrJFFM65rbVrSBhwwt3POeMuajBtzgrFAK6doqKHM7dsmXz
VhjmMrJ/U74uCx1yXW43VBJylQ/i+YPRgKIaATqpZ4djZjhq0P4xmfWewUEI7p8BarFg0jl23EKL
rk95+wlylYiDulI0r9dYN+8b3gdzE1x82+njGf30ekw8blWztxH44A8fEuXjNcgk0Ot/zFrsmknL
CABaX+qREL3q8N7LSCFy3olJx1/mS1VlqykZqpSu90J1Fkz+sEGfPGfFHKlwRPi33/BXL6O9B+NB
B89VyYDEnN8Hhg/eFM31CQrmpafnZeUikzC3rtTtVRSjzLTdBKgZcC8wSOGSlNkHOSbHz4HQzOJu
vcG8E+SJvqt9NR4bIoZABH/aSDdmZRW6lVka/thALzAHp0HH4JvySD8i7E6uAsFwOSsc9D6Ik9r+
vtqLy9bGS8QUUixF+DVeSfyxqDWgJCHk8p+qUtsZZCaMUErsT8mnA20ZmxIBEXxy7sTqe21bg8HJ
ChYSnIMQJRP5LBTUVDX1pcVnF5G/XyRYZDROVknqVxWieS9HvFXmTsJmNOz/7vdLUAuySMPf3Drf
Fm+AtvbP4tzV2HNrg2VTYJsP6aOWq+BAD0XdUpqaCc4B4qocsCFvY9xCXah9uBdkmxRhtZFlvTLv
Ur7LOEjo1tX0d2zMf51uuMBRRjJM9oah/hXwfVqtArPXq/9WZPv/itYd8Ddk826nH1L4R+8puQ5D
+RoZhNWQiC9uo9KIJ1O0O9W+V98/fYArbLqEU6MfaYBVyADmUt0Fl5ks0Jdp5NEF2EOHf6oNVP4T
ARcyWfndvoQmIeja3MoUASlQ+U2tZbqsUSak43f3VK5Z9WhFo0O9cGa+Aa1JpXX87+U5DhJHjW1k
7T/NSFsOl6Ktvh7S/WrBBJai2Ks0jwwlR6r4F03Fc7Y1RsNzEej7rXy8uGKl0KYl9yAbhyJpo3Mc
v7kFtKp6MdUVDk+PSQDMfb1E7J44UHoqyJwgl8Jp0mjdSgk+4rrJxhagzJ26l3Uz7E9EDt2wBm+2
O555OZjTLubKBLSMFgUcNrC2qrJO6w5Z2eF9lOfWjl2tKhPI1m2oinAikrJCLGeFty2FFi8eG37p
TOPTCzGSrtRW7qUoJDwC4EizqhlUDu/mGApdjZyKMv28nr2plZPXNER6eUFitTWO97ofoRe0u0Oq
ful0V+5ZxGKld7mRnU80R3cV0y4m9BgiFV4RDH1P016jNCrSWDAnajIHqQR0vSRukrjn/z0JCVOU
dbaatpndjRQc0mrkudUoysXFSrv9OHkkC/lKSzxMHT2FB5XqQUz6tKY3tB45Se8O7fKfznxt6+L6
QawHmuw9ux8zlx6sF20vLUL0b2ymyfZt4wAJ7/1BC3E7IKaq1PKRK4ed4+8DcboQe1EsKcT7YWcU
ECTE1i8c59ftBnF+MwfPngJgoKGBsPiM35fcHHfMjV/YKubwK4lGCECGzR598EbbF8oo6aWPA017
hf4sqzhJw06qWDVa21QjUSz41RSAsdrYXT0ULbmuSbiY1mbQ+SngynvIJRNtImycC2F5u2r07wbq
ywmU6V1WVF+PzCfFcujYUtd3hioyaByAzzjY4O3dLlEjUzbkLHEwxLgmvThXVOmFqA3hM5G65Jyz
zAk0wWsjvlD+nyG1JgAbMTVQn0+sZzR0t4Ta1xPnPLKBPiz5MqXu4QBOt2dwpgKOB9xmhZh0vSry
bo/TZoMRLGkZC1fyh/Bny9Gb5UubL+7DazQejVCLNEf8CimYct9UrK2e8DXuCzgWTN4a4iww3erZ
PWcvT8QIT0i1E0wPNt8UQ9Kwk3tTepzy4Z69IMnxIWQFQntZJ0u7eO49Z6q5bgXE/Flwr4t9ZnRa
gak3pDkbTzxn3l8yLSSLv62+deEUwMzFyXfkwvOH9mO8gFp7P5N+oRX/KsMO9QmMsLnrPaNO04kh
UrxJO2lVTRhh66womdZ4fRIDFWKKkfPcR2A8K4yKcPH8oeYHysL9FC9Xkwiv9n7++6/2DYoER2zq
9tZSItNz3cOFZ8HiKpuCWEtUZnL0dQ2DhAOc2h26KE+99DvCwxgnmRHn0+nfUCccUH4lbHGZqsTz
Ds/5yhSVpXRKByZeiaL0PUd/Fa4BoEsZMj3MdmMVWlMNUOsoP6/d2CwuQm/DXFLa4vOjteVIkIxl
+0sCmloc97+2N89tEFaycDLyHfyWi1ZjMtKoZZaNohH4hqcTLtE0DokdCJxQf74OQY3FC5hAI7E5
n7Gdjqmii3xytHew1mk+ejZbSQdjQFQGCO450h9jFWsZo9qy+JyaVhrNifBSr1mrR1SudXtz6T6v
wi4Hz0+WIkbM+N4hbT+4cRm8tgRSiptP/G/aSjyVEwYm1Frjjs/edMtbUZ8oZENIiM8mIvApDhHb
ioHFnNtqCaDJg3GrImVs12vejzhuOLNICFVtTbE7QEfGj5PuvTfSG8TT5ED41q7uZ5fs4/7BJeMB
rit3/xhSf3yhGIJL/U4ZkPNeks2PZqWmVF6XKQ6pBnGEozTl55QPlThfSeHUQ9I2JZM/NbNzyZLV
gGBTF3gcA9Gvl4NtNCes6Jk8avdJE//mCya3sfJVDQxgUUHqT044JIgoK7xPH3iJbGIAMNrCeSXN
PmtfeR4nT83GlqvNnn8K2LgXjjkSsYWfM+gp5N1sPOMyt2JNpxnyJsoABU2D1qegBLXD2J1q4VPG
xkBXJ363fkzqzyLd+Qs+L6YUknfnsCJJNrM57ZZiUq8Whiz+WK23+q/H6ZA2Icwd1MCJr4kmzS0c
qlB7Q/nDAVqlEhSI7hW85IW15IwlIS1mkhwKKBVWbz0AO3mTeXCWItk7WOmuaul5XE1/HOhSD4oF
d5ha2ODI3oFGVp6lbS195iGO3Ok8fyE1BGyyoP0Lf3XuLrkZuGBWcY3MfJdHik52TBVy7ErecPp/
Hu/JA46Q9vpwNw+vH71u+NYQ26iimvdLOvOZmCxCOmlkerT8GxKEhNCeJh4EWd77Vqk1MOZ+W9i4
f4y2kM/D+h9+UY7OKyaaxSR0A85sUarB8E4AkGGBUxds72b9oYpBFnRHPRZXbiyUZteN69FtBO52
dI+5PKj4nUSv1p1U8Nd9a8dSJqXL5Z/aUmstt58fAWTkKift+guyV5zk46oWI0n+qrCqI5kCRZQ+
SH16ZOk8YzByoY6pU8kXSskIT2r9a8Rjzc04jv5Du+APeXsMm1qPaxCQKBviFzISdntzfw83hxaM
MY6skYVcGP8gzqnLX9wl2ANtcQCs6h3V99qWMOYr+uwBFJKiAQOpT9yepkzH9VXYk3aLNjYGlZPR
FAEOalENGi4l6Bv4aQfP1kj/EtRsq6diM+GGs/6adl2ACBI0VDPGpMxobngAaWH8toqaUWstZdSU
7XovDOQsdtSktdTqdBfNwiXxaftjkVhhtKIdALtAP6Ir1zkYpGMXWhJQFkTB2XpT1uOGnR+T69sL
8FLaOH3aw49wlmu1ujnrNbHWRPRYL/TWOHzorMxg0hhApEqCnYHFWXT2VtS9rCoRqZbz1iRJLGVv
1t3/jF0UgKw1Rb6DuX259y21uk32mR6koZkOrj/ymu0Qc+U9jVwdOoVa8Glq/1UuLjkXre1Cn9Ju
FlPQmoACoZ1G51AyruRrqO0gZ6QyYPd9MUoiQRcWoxdRYNDw+wCyEbu3zRd71Tw+55dfW+1LG66C
K6sKcB+tlpe8cmsQ0RJ8npMJgFaUD7RuhA/DwDlBywSbgnlI0bEUrRAThzboPItGHcmFnfItuyk2
wRuYxUajyIfLVJUSbgd2zTUDi1q665CMM5UtaDhqF1nykaOnv7mfD5x3mnyejv5EyVqd2YXH5FcF
YqvNlcHOkfWffMyB1reZZma/qT4FghMTveJWb9k2Wur5JtNSuXLZ6yIHkrkORlIQ3LtH/MAHmuV5
v9eYeC4RUL9bSLxYxV1fjmQeN7Nc6Wr5+8ZWeFwwJkAZGF6CvS+iQLrK1slMUewQVxB/zGEiM3ss
2Sno2HU5+OS7jCuc9yra/qPLs6OWXHZuBKQl8BPiv4tuqQk+nOcuAHpdc8oMYGdKlzCl/r6wIXfi
67lUFRcZTcr969IMng4t4aBpCXTEzVImn1oBa2v1tJEk+KfxKEeU3EJhCHcBrNGfy+Sw4TCGcrVW
1nMsuLVeOGIRCwnP0l6DvPGBmQJnloyiNyKb3djWIyzM6Qg0rvDMIcFL8gFsYpQpHsuHP6g3YM6y
5ZNWSPqRx7eV7a0UbRQWYq3VNviPdvJszMCKIhJYD1kq1Drhr3RZq7f3poKJhxocqSay2VKkQCGO
K1BuT5KEYpDh6BZILhzoNld7zfF7vUQX6J/JoC2FCeD2kcETY2ruapV8QiCb+A920myysYvgVyU2
Rys+syZ+dnRA9U27MpS9NgMLbe+JAicKPlN7r6v7lHtG/+pt1GdMHBuCPwrR3Wpe7GIOxCLkkmZu
Azd/9JkNvs6wPq+MchJIgGQcIS605rGpPwOCBw+q+9q5tLMQrFcxcIfoh+fHggcPJ0xv9IXpTcU8
nz2e+k/S4fW04WXVRkG8iUgtg85KXXCsk9maDdSXbaZnxOg4n6Nx8xW6JTi3zbkzHQUUGLhWSgEl
G1q9gibVFLhC4HCYLP9J1o4R0gNZPXS045Yybi0UY2ChkPu7vGqilkQ7oKpZiDpN4zkafuyai4us
AehommYGgmTe4MqC4pR5z3uw6TEKVpWUGZop9p3KhzUzwSTztLDKx9/9YgTNfdwPuXJPz8rmTQAY
sw47MZ8VwD09ZRCEL6NQ319PbSAkeB31/DkYb3YMcUmp2vibW8Qv/m8/hkWhDlZv78uLusj1kCTV
p6a8JqHk7i188nWLMabxmXNSgij4Xn2UqV8DVnBdoJk4OxrCOEQzymYOwk2BPsVN7/1eqr0cAXU+
jcJS3bM/Mx4rcHLnqg4m7iwBf+EbZTRd7ohGmK+zRsW6DU0ZulQHJsp2YmPoqCuyRo5kjMWDq6Gc
pcwOq2iHqTIVMdlZQ4v4VAedwFBKie0KmGJ6ji8YFkrAwyt8aFCOMfnmwkWL7sFifi4lIoqWydsC
t5L32l2oZMiS3uf+fUK27DBsdYtT2+ZPsVXeSEUpnk2YeqmowlbJ9r8/ULp9/wWEKSipORZcwnwD
Nl1VxCNv/Q04JNjmYvx/X9VjRNGUb5MzuHfZ7ddzBBnM6m7eRX7D15uYw/bfT3rhUKaGLjbXuMSK
quEIez4C6sPcW9EAR6DQMxdzb6Sy41G6KzRxQKvtMiYOkYag0b+HgQ2MOApSPzLOgBhSrWl4bPK6
yTM9X2Y+kJSfFe3mF2FrbG/GFnTgpqLQuS314HWKxBcDFP1pBkdLFvHiDBs2acn5wTedhwlYAdhD
mOivHi4AcwDGWBdr0GUq+VwiSP7Jv7ZHbiOrTH/Jlsazjy6KIrWWdo2C1/2nVhn0KIAJE1Yjb2q0
NGlgluWiWJZfegCvsKoVuM0kjsddGwzcavk44wpm9gO3YjhlCl00yogVit7SYKgiHARmAIDRgJ7H
cGb3TuIDReGVadfX8UE176k+SvBlylzuLuSo/fqYjoSJNgALwXoU+O0apVS1MTlSANjovTOtoLBt
/S1G0xXmKJMyNbMe1qroxWv93g9MjObB5x2PsVicRXFzSLv8qK5l59/ngDpcKSdo0ARLtzVUsZPE
vi0bcxg0nypADYw+c66PJzt7LOjt7A9yt7/7jBSh2t/h1yhu09YUrHuGJzj9RY+GzpLdaNqRo+pL
O7evM+XfBOfXnYTIjU1HTV2oldgrWRbgRHJYwN4qvn5PVwrFMQeiydaAdYOGdH0iVyqMZlsAcghp
HCEp2w7RZsa1fKYi/fclxAXlC5MS1T6Pg5hDPVnk8EMBtRBrOLeXlWA9HvhEMwOhM8EWrcH/3Qlg
yoz4HojFiNFeavjOsQ0Ob+65yomH3jbE/Lv7uaOc1Z8foZ3R4KZ5i+rNHKbJFEzGMXqxmUEFqJUj
B7NkKy/vOJq0MIb+ozGdsKeYARsgWWOGY8EqrFEToJ1c5GLikXfvAVGR0/DUfzMGC1Mv0LgXATv5
9F70c8zKi2iuvKydKRBvMY6O8AjIAIt0Z4nkj1IPT//AuDXcA0wHh1fYRjyKHkmGqtbyCN/AX1+W
ZmJtdzyj2J8DGV1IfS7gwRihSj/KlhtzBzhFrXG3ANfPkCM2RcZYY0iMv1jL8RL7oiaupMAZaDWJ
oZk8jsoQ4GcnYZZxsEBHShltBcbYuJ0ygi7K7kgmap/JoDupolkGEscc81tQ2hAtgjWrIZevDVjm
P3qEPjR3S6tIGANhRdD7Kv+odo3BMjsVSGEk0MPYGS0EFepjFFckIfbJa0XUjKvV7vGtOkZME9lO
hA9UI2GRQMcPaE63in4NrcK3BV5FKIzSpB21ksnkDy/HXs7MOEIhrVkLrvY2LdSKbAeZLanhIdQc
fmoXNJJyaCbwQ2RQVS0mUfo1qlv1q6ru1Ivz4WzKrBKMPaYxkwP12KUjRJEuzQAWJuZCyRkPu1ll
tViwl6NxvL+KqxdSN4ZzQ5Yz9AnhCSLzEsBEWlQDyF+5Uc1VDhTit8Ad6WHlgM166gyVhr5N+n5h
nXuVPbKm2LW/k7ct4eNAMJsLcg0eDV3LKkORYjMkPioBUrqwPAJr5be4uWzy+KjeYlwbShWhatSx
33v7rWtn/oJ0zp8oXDtLP+Y8cj8c5f6wt4mAwJhxXOyIvN4iuuKf3ae4ElqrD6ZQ5xUKpoUOD/ij
gIJM1RuNaj4pUkM/UixuBL1whHPHNuWJ2YI25XGBBX6Qa7t86qi9N8fpbdiQmWnncsvTcaNKCOcZ
gjGp8kU2WOX5o14TmupQ0wgAU4oYWcinRRjTSs94oUnZJ/+lf4leBVk2HmlL7CyYeOXiwu2oQLgv
fYvUiFEHu7KwKP8Tm3+OhOGhPE8ZZlkphe2GoY5/Lj4poSKCccUarhU9qWnn78TCXyxza5jYkIBE
y2MjYljVmI+z6ItgUtBqVWDJ6wXXZOWR/za50mwCaQf3yaDWUjw6hDZfDE1SoXzmOB4aI0Bharnb
ustps0EX0QoSX46j0D8LvVly10mfggTUHykYpGQM2CSEUacfkJCynedkUW55e7Ap3r+h5G2s1L1J
l/erXrL3jbAH+mB+2bcj3/s0y0ugfccAZaKWkZBnrKpL38MkgpN+HMElgzv9etSIU5vBpTDL7wqu
lVRvXZE5N+ICJEbCxncjXrkpikJNWMx0uODWwBX5j5LhC+bqBlr6bCZBAdtbhviJnbOencGGMDh/
PP+Ji9dG9nVA1Vgtjy2xk4lhfHD8wDKCx9EDDlY2y+6Uypn+4PKb1TCY5oMtsqZVjZK0FRynR6B8
NJa+HI7GWi/iBdEtRF+HD1YbRO09bhI+P6/bgZj4d27R/tc2VEiMkgv4CSmtWi2ZUj9q1v57z3J9
YDKS5CQun8jmCg8A0668YXGig3pL1nP5BhuqxhnJzKobcNILkTnBqkmJrfk3T5C8NPdsDvCwy3a9
8NJnpDxSqPnc+qJMYOFo04JDnvjaK0woA8g++2LliNxkW2znWByl0Oq7ZinMlyQMHbgzZU585eGF
ZIBoc8KFaaEY83B5Mf8iUv6Z2fP3RlOJznw5uDVHbSukeWJjrdam8PUVgyiwKD7C6vCDJ7w187t+
z7iic4yjIokrjPrpRpchvqQ594CDwu3mxHlbgsjL1K7V81bs5DBAoDKZD0N3TU+vq7+Sg95c3ieY
edbgJSnVKS4JJ6I0vWryBlzKscA7PIS3wBkpOUMSBhDGErBg6JxY+Qnwaf0gmUfQmznpG3NY1w3g
vQ9I+nTKuuBFrS/qf8TUCWQ63Xjm6dUadAxo/7R2tcu18hsu5Q/bkO8QsFRUBQK4a4zSMbjmw1Vt
cNqch60HqwE8yyaDPdGWNus331OpGXmNiFMNIadFReoarQtZqNFHWr349oNfbt6kB4YumpLaysBI
tg6r79JOOZ1TdZEhjlwHVmbqa7QDYqtTp11qtcxwuNwaOJXIYewC4GTeYf5YBbCP3Yc2CmW+8Ted
HKQORsWO200z/4dHaM1/eyrG1eB7ugo+cWyEWEuBOLHKFF6wgWNWq0TpLiuol/VsDZ7QRGgz993z
yDRxhCZVUs1TCKbyxh7JgD5zMeJ4b34chdX6Ykk88NHGWz4P7+NNUcGGaL0bHUhcnEhm1fjScTfq
fN7f/kWPqa+7auBNOS7UUrWRNwBEmIo9WT7UiICNIrNeLW5CzYONMaz5V/1hYVdtxck/rYyEBGaw
4HvY2X4o1VQhdKfIUyEP/PaIDTatcNAb8WSvto/bIPl+iaCzi5pLRiH1aGSifKRawfINQFU15SUK
w9m3349NmztsG0X2ahsA+yFCsRqAqBTVgS/rq3CTq5WqQuxjaYCRGtI79zkBp5Rtk3uye/1y9AMW
qLG8GnpnRbfn2jf3LhJ9i1mtgbeX0vbCVPWSDgaTnXQk2UvgRuz8O+JwRMQH46CkNhESbUAHMwen
H1hcbY4nzV1XCwBOUffODS1V8PundQ8aZPmEk4oYJgr8U8V3+yescsv7T03MW8IEeB8SRqMmGAs3
KrBlmCDiLM/o72l+7b65hzS/LWDOUcZ8j9RSCuf/32m1KBJRLuMf4bs7OJajCH2semE4lxglMKbc
q8XVdTa3Bx5oPSVPB7ft7MtZYTYj8rdu93Qh0sO5CyQpaTMt8Tr0Undbsa4r6mT8zBxcfclZFsqX
ci6uU39C0/MNRpCHcBk7sVsm4fg9klbrkw3zhe2fJwMhV2YuaG5jTl+VpuReIvJYPLAP388MKiNb
BXxtNqc83aZgt5+8bDEeurfwED9BDq7NBL4w3j3eQ8FuS7N6TbRk+HGMfhXI9Y94mxNFHJbbEBDU
KRDpwovQ20KKMmor4w5fMROwQ3WNFBcCasDzbhyxeUE7owWFEGoEl86CnQMWe5QbYDJrRVnazRZC
GvMaqcrOwYFVQE2NoMu93Z3qWCLQ1betBq/ezNnYvqCIGboa1WAVYXmosFA3/wEZaxOIPtaPdriU
aFswUwH/JysSg0oE+F2I3Ncp4RfiVVZuMlOIcSnRU0DMj4EMdvavQRVIYnkS+UBQGcuOLKC9yawx
Ez3vUnwJs0yv/KKqBIYQJ9twdzGZAWPqVf0CC+IcOPOF4RZs5tRBt1KQn8elcjpTMPhc6gjdVJkz
qB3VOurud+qhahafqSlcZLmKv6GVGFrWyWVJ0yyzTCN8la0L/vJ0/x/salSwFphKS1sc+nhB6pbk
HtdrrDFclznCdZnCDD1xDtbFXtwEzGVIOgtkED5cIxNWAW/CAFBx1EXDCcSD4V86cpLfZRhgaoX9
JPi8KwbXTupIizNJQqiH2rZJ/xSd2NtIGdt1vA5Gutwltk8PmZjQ8ZrNLEB/DegsVNT4kYTuLi98
PxWdeBTG8NFXMgGNvsa6x3zelZ2CSf2C+8MfQ5lYEVl6xRFedxLpfCCk0mfcXrDHl1JaipChkuhF
8+Bb4DOkqJtf2bEZVD/IM5cvhe1varceHGh79lVCdtcrRwAXQqauK3x2AJfZGedj9fTcIgwXF2B3
qqclrFjiCqPcMT21JSioPkH3O6c67wxeN/M6J5+BrpHNjRGOCyiLHhQ34l2P9Og3JhZJb5su7Q2v
xuUs1y6Ouf9hqZZcCTYI6uFABHHcFJtUcInjFw8EU1orb3cBaGRc0E76/sa9Y1H9ihDSU4qQk+Ck
u787LnLK1RKhH5+wGMOh27AxtzuWd6fAg3be5OtcYVRvQCn+dY1/p51qOqECoR9iuFuzz1u5r9Av
4u9Qh7Ck3SVldZ5e80FM8Cw008fd/4PTQ3eqT4/QKyviZdb+VVxDgZP3B8533d/XSHitq1bStw79
ODMCfb3JkIHmBFOm7AY27rdi1eucxUPw/LTg9086bi00rvf0iPwlqphRitxAnDwoQGnX1UVe4RDU
e//zuIsBIfp2lL4Bt4jg3J3iiFmNncTGs1QKGffjbzBbrlwJ7Qgckm7UPBn1EA8Jl9FsoCd4but0
y/sFgESTOFeebC6lciILZGah/YJzuBx8OU8NllkGAh4mypma38TN4Ti+qiUOV7bTtlOuC/jEJOLf
TqC10bXk0Fq7dOErQpd36lReA1x4XWX0j566zN9wUm96Cbkxf63Kdr5bZ/k4oiZyUsP0aGCnO4MD
Jg9H4461x9xLtMoO5+WhPQe6iaAY6ckGqxa8xcQ/AH8iEP65O7nziHH8rqHc/UDTR/e/rlLslO8K
WWfvpmKDFt3TkvNMSKnzjzkjCcTKfQBZQewzqVy437G7958dyQJjtWgv0vlOqvf2YU0Xw9bVsRcY
wiWYUJQz18lpvPRaKc07dD1/lhshG2K5hq/LBb+qWt4rENyvT7PIBD0394AEOY6SuCyQJ/feHNoA
/KDVdBSuYEhjirzJiuv66nvJGDH1lQ4TD91NuBlUFCo6rbYcRU8m0kLeAwgc3P7dGzDSeCknZdyr
PANOpU/TSseebTQLUdjE0bet6rGQcVTp4jDJDuCUpEVWtb2z41Ak3PSrZrbmqzj91bUJvN0qO0Dt
SzlPnYQPlRdNEvfZLM0h/1r62RydptwD/H/6CcQNDV4mP2bld36bLSFvSN4jYIhsoLr/cq3Lnjwk
a8yym6Wl1w0+pI9Z7f5x9HtZx8LMU6NEDeuG2KFEy9gnw2xVSbMOyq4n7gVuYvKukhM5CV40V60s
Toni/bgdYUiFt4WnVc/NpoVRMQg0ySfv7GXhHYKDn054mHc2uFJCxHAucV/k1tp0+MUr27IDwvGL
5lrHZlM36fEgnurmy6/vL88+ZjZ9PO+hp4VONcyIiBOznuhjdbIRfPo4x41UYVRxh/hwkOQATi5p
EtBTBtotHG+WFPLTr+Fna/qM31q9WFS05+w8m5/Z3N+iIyZXqwRIaqZ3SQo9oEHYaXbb1ZVBBZ//
m2U+M8dBDYeA4TN0jaHIsWlOvckNALED3oYc3jM5mZemqDMHfPKq3herGRZiUNokLpqVPjiIjCHV
sIIdx61NHDrftg3QOGS7Pfc+eEDCuggK7zsHwGT3ujzxgTB0byxPcgrzz9stq1MGYoJeDVTb2oNY
MJybAjnW1zdAST/dJOSjsISfjyuxiYM505pz/PzVCZFt4uy3dxhr1OILiaCIFYD6KWSW6VmHiXfu
NfpL97pIRI5uOxZy4hwaZgJTr380OYPUNOJgGHjys6PxbUe2iJIZYl/StFAU5x0lwTqUR/lPOves
CoWxL2jFGtz15JAzFnZjP16pwrsxq5qKv7Ucbi3ovK4+lSPDZIe+kK7d+0NwTbHqbFIN2ImPRySt
NOQr9+2PtznkjabMM2a415dhITAyR2MAYEGy7WnNxIwKEIjVIzxi3cgqHIVwtMliQDUjwmq6Pirb
KYD+FDfhiOrn/5x1ximUAeY9Z/Cqi6ljiRVBX1sDX7PS5YvaY/NNG5Pvjt3klcbRCifOOahBE2gX
5yQhISwwg/UysvJt7HRScjPey2xbGeVp5AXbsjBw/Dpyew7q9pKCVs8Nz0gKQA++ifXFjludeSAd
gdODYX37/jYFtgPV74D2aRejAdzXEicUGV6u5hg6UPMbDPlZcHvZjh1w9evoggswQmjRMlzz4ocU
TYxODVyACCC/xxLRLKJsPM3l/Js8tsHMSH2y1z30BjqrdPZwlPTCYslGzbe3PRUifgIPhHY+qzqp
I6N2H+z1zovXuxsTWV1JxGO9JfhWWxsweDYP36Zls5Zb6A320r8OIdPbzFug3uhIsJW/5uX81s9u
KKQ9FG/R/ti1JfXGXDg5SZ0rSuKVxujgCas/RU/XWm7i/3R72egYXqR2Ss/6W9FSbxMzth+FpCgm
+7vqHcA77+pXXYpM/vedOnKZempaWiadS27oM1gaQfdQJQKMoMh9zUoIeietsP5fL8xSO8l3L30h
E9bfns/PaV/7WBC5N8qcjtUXFPy0ia/FjNjtuYVm0I+0Io+LzPY06TNH1nQS6ouE1ZnH8f862DQE
z2Lc4VfTg9aRxz7BfmMNYlvjujEV8v4ITSmSIzHLakHvm7jqHssJOWw0gFCJs2CQFYtifnDNzm98
i9z8bS9FL+0dpI4p4EMH2qer6lqFIhG8fZcTTB1zRbRLsgUbsr9+9uFZwxFWLupopvUPwHw3oEaW
NNenis9mU6Gk3HGwa186smJ17UEb8ZO7zKod+9leEn/mMLl1YLaVrfsCktvAH682KOZw8tRi24TH
vNA01VMe2T3YxVAhvSf9dWougqB4KetXpCLYdHlGcd0RiDGkGvY1kYVMr8a9ZW6C8MBGCkdkTOK7
JUs3PGhTfZKSKbovBXa+9u5SlQ8gccb+5Z6R6Ub8bDcY0XWaSCIE9hm2eY8fTBIIBEruaC8a/hyI
dfJNh1jFhNzuQVmoPONjgZX0qXFDSlDNfVuMDPL2dviIocACDJATzyPZZ7jBnAueKAmqq6lrDwT7
oIx+X57bvAbdeuxTmkxYm8P5DohBnuxJptuARlwWa5N9YgAN+FaQZDJBvC/IlFkzIhlxfCVfAb/i
NKsxzLp89z6IqXu6nXBb9hzJW6dEQS2rJSq/r5J1LZlRCZzZXBaow+rdBsQn5+M8CdFF1ogotrJ1
LFGWk8Wi77HpfDc/iBw0K7VRSYcmoJb6wcm2TwhzyA0VNnr2gFzeIKlKjfcJv4sVrhopAygk5Lj/
4NUmZr70j9zU7Mb3MjfoetEC1+ruunHW8KgHKxFLfCdWfG1zSoLb81vBmcQUXwaf/7/Sso2Wb9r6
qhTNUv/0gfn4p8GJgk99SC1EvFSl7sk6CqmiY5+3QCbWVPsKHsjkQOomXVDKISr4/3gtgBIPFYW0
hajV7rc4xZ32mvZy/z+wg5ztMhKM9XjuFdX0IGXsM3Pk4J8nPtt/Mq8MSWfdw5t5AajZDCGRuGlf
SmvoEiqhaEZhRbkNrK0utcCOtsVa6Oq00lr7AQOW8TVzrJ4XVLo1SfFn0PlIvgeOWVSZBfgJTcby
vRW3cdYUghtbWhRY7ocnrfb7LP3et06+Pp3hsuQUQlicEg7r4v+DqLnJf8bN8uHNqDdhmgazUEbA
Uyj3NZCEFMviCrqjoDldRargrCcpXat4Lq31NhW63ee3Zv1NM0/6WhYdDZgCLKSC4I1OZqKItpaj
l56v8lIzHsPBHVMsQP48rI0YAqcHeomq2mw65IqaC/fMn6OaBLE1mpAkI1Iql2HxmFdiOzlr/bYw
dcKLdWh98OhTZhRusGhHWjldm0loI36AAyt/7oD5QVQxrGq5LHNUA3V+dXYL+PxyskOTW7PGpTui
EiGn3YeotXf7WQ6rhnJ8droJX6fNc0FdQ+wFtR2+RDpgz9vrw2o3gth+IYIQ52Dkr3obP2A2P4w8
EUEK4/WGLnQe5xnPzIX6G2KB85wzvDR2deqWi8oddvw/bRMkNM7sPg9uzw0lspiQTFkq0wiAQiC6
CzItRTQqZxhovBk77K9CNfcePFOca+VlwGmQZq7blHGLkRbzXcQ0yy/Ab3WVlHpHDyaUrWJLmpTc
/V9C/iFCY487g+XUi88QgiWpxqKObaWmc4HOmPrltXQwg8qAIJ5OPNY/RoOiCpxjw5wpw6EvCiJp
r+i4BMburWlTOqDmZVNP1xr7W8cGTI+jmCzv4NP54+u9giinhSYN9kBlx4CMnFyYl+InhF79xXBe
bAxgvhpE5ViGYPB/8SatMqPGwfjFZE44HKEDzUJOO/6m8CC8ZrmE8sP/aYemRXeESOBJGVylelGY
gVONBeSynepfjkXtFl+P9CVdd//6Z7PVN0eDgvJ88xkTtsJb1ZDMxxziVjgT+aD8MI/4GhOKYl57
F2xS3BipBaD8nEPPXXuW+xOg/FrcJc4rG5X9mYP5dy3g0sZz9o+HrlhT5hcOFvxYAS2HXgGyRr4h
Maa/usstr3vs9PcG8kBGtwPRlOthWD9XKKN6BuZrDllomVuxtcMNKu9SqAGr5IliN5X2K9+oD9UE
M2XLN7e/7z7wQCdz74TNiJAKCLwdralrS1YuheXjusqoPcpU00E/RmlvrODgQFd4/LLtOZGs9lmp
Lhwk1AMGWfeLQNuHkyt3fsDG5CD/gyvtrY/BD9sS+kUq+WquCxA11g8nA9ul8biQU1aXv2reg8mw
0uP1dHkN1/2ePtThIoMLiX/d/WEg5q+QHihSvCVN/IPBEsC78t3hgx/iMdIedxgK+lr7D8qRZTam
jgbLx0slcyHVvgjTYxrlQ5bhsX5rJCJADXN77XyI/FBgNBXtg7KsiPY0LZzOpjU7tQdiESkpepMr
RTQUWl+taxgYUDh8I5DamU9n3SkhWIhTwjWX/VEV8+onX60DyrQs4Q5wecB4a7bcZVe2cJ36H/qR
outZLZvZgS/uDIDVCMpUfMd6+P/d8gZtB7uIK1RVGh94zn9ZD7Oln/TCZ5BebC1EXP7zGpWZGwE0
hAQ9aK/A4QcU+bp/j/MpuKDPzhi7mhHCbfnNd2yYCkl7HUmV1Nv3qjeVNv5PyMZ/eQIkAu4AAWI4
ycPIkoM9ksCWYxqiC3vcrRGDSJE6fSaWAj2ET39gn0Kz/bJfKgqIxuIvuCNJ8L0vsOkogRXMbu8B
TQPJ9bViIYpuQDPIEU5Q5cP7ky3VAhtxlFO/r4ff+hRK+pwnV9abn42N0k1zRwxXd1UES+IzGN0T
Rpe40cjyp52ByoRPye3TzZi+5r0FLm+Uw6amLNmggaR8jDm1qgKub0spouLYPKwfjiE1bybaXjfB
ElMOyx1pTWCcoQn5/XPrRSvdrSLfsbrM0fegTVhrCMauR/wbDyGRqgjsbYQ+cbJdkLAjqI62FtA/
mV2JPT/nVc/vvsNSM/JzAac4uLRdUSm/Yibg0926v/qoxIVnV/0G40GqCCNbtH6fiQxzgitT5nVo
2ISB5dKNPqi1Pvv3kAg5oPtfyPY0hQ4CyU/GZxE+lXHW57eh3AuqlnbZSLDPROcKmFeDq05drI0V
NEmOCgdmxLlYcSux1mqjiMFwG0Z8XX3IQEsUkEjrmvLL9NvxHLm52yzKVWLQQze9qySzQhcQsVfy
a73UsmI+8mbetRm8Pj0w0M58S+tI8cJVyyfkt9/Gop5jCDN697ulHdxirBlZ+YWHcOwnDNRiidXk
60hLaA7JPgKeR1G0fFK1HjumXlFFnGCKIWqGaG0ssY/Ew+9g1gFqYRaE+sISq0WlLZ9ZRkPKcTdc
i+WgClL6y3he9ajjNetlrXpDR8jnYg7Dl02ydclnmcmlslU2G8vXPvjWvVxqb6xD+xWRuM20yrnk
1jFC+GTdfwN0Q1B8S990ObIM4fiViAdV9R20rdSqCXtPbFjRO23sX3BWiPeyJOoQcToIQ3hFMBWd
Rg/SN8EcVv5jPtRDJbVz/4Hg5znTPXsBAxVjYXqU6weyZQyvxjISCkzotZuEMezHUxbFcK7s1StF
6iuqWuUSJxKS+bxqPdXlksZkB+fgYhENL+afeaT3EHasLA3pDDJllABGsIB3Y+cZcc+GkdNHmvc6
htHvg18X6bY41ZFsIgSXl6xZ6jJU0sM0MECUUJ7fzTjdcw1vZvFptN26gK1WddhaNl7TDgqA70D9
1nE4OY3On0KjwSvHNFh8jzYawp0YOwmFePZYmXkucHeM4+nJLUtMficXD5JCePDIMiaPeHvowl/d
U0oU8HMbTdN9EVpwDFplgmC1PbI9Cb5sSGM9P3z2pabQT9nLDYZUzEDs1bFgS0ufi2aSfyzIKz5Y
wo5WPaMEmoiGKs+yjEHam2I0ItCJXYHOw40VMgDWA0YwS8Nd+WkmFB59aFJZeI0/r/SGeTt7xM0S
7xDINSfVTQ1qy55f0l0dyRbxIerqZDFU6pf8Q9HLYFQRMiL0thJh6lU6seg5baAUxvrB7Dh2Tb9G
T11vElmGB0y4Q6iHKdQXBvYz1Vcw0Vbj1JHFA0HkkLjTEi3CNWU+n/pelhGwLF+sGNrtxs4PuU4V
oaenT5V3CQovSozBoinuGsaPFr2eGi/Bo1JLITyd9h2EbkEzDkOIOOXfE3BbV1+pHxvQg4ohYMME
LwWu3D5VWU9whcdmoA+OKChbEfNkTT84x9rxflZroWSqbiC9fBWRZdPKFies95cGhnyCohK2vrR2
P5wEZhI10i9C+BHYeCDy4PrTU5xl3ioYd6cEZgqHZHMOrOzwM8oRYDRlbMQZysjJps2ZZf8sl9fX
42kcs3pxhEFxgfJhDD3WcBO6cPmrTi5yw9FSGj9KkO/pmWRtK4eKcSciK7Icpdvzn5EguMGNxx0z
/kjtexz9Qa3j/boBq7ooc6S+D2LHoI3uLlDFPXkrPDVTiPBxgSx/H4PVIDRvIcSgQGROCV/ZwNkq
cCLlrAaLDYkzGCAjrh69Fq/FGMXm9BKwE2YRJDKxAkkqMgJB9sLvRGdglQAuZ8BZFwNK9Y+bjwQI
TkLZAFIcTBMVBcG+EtO8bIUxS5cx1IWyvV3pH+QEOND6UZA5gh78QuSpynXaIfO6WQ13U9h2BR+S
fEtvAOa6tRxwoSREfOzd5tziZhqf7VGtRIZ3t34uVAwdbFU583Wig1FjHkCaoz9NsqlIHz6Vne9W
Yof5P4VEvOuLV7llyc94sw6dme1WEEEVQsTIJARdXVn8x9+lGm3Biq+Y/YtSJk9in70vOKjtc0Ir
9mvAYcGmKTDagWbiMq8nUhsLMlM0MS0mKc5z2aB1Qk8ejyoD/KkZZotKJeqP3JUoSgIgNXLLxoOX
gFr4mzK8XxtelKPXp4QuD067oq+6qLXjmpu37UP9tPDKl4nWR+spMyVk3teMecmYQ3Z+RYQk5j6h
1vaJCgtO0He2jTjcE8Elv0o9hdMlgpRcmpihnK8rPjIXpoRc8f+s9AGk9rAUhz7pcG2gKsHXHDzE
DgY+wltR2m9U5+KwkL2TI0zvKcxhiMTaCcSfw9u4gScDCVzkEoPjUXwjAa5h/Ki2Q9EMJn2uiicP
M7xyqkmHSJsfyYLW7E85miZHtEqy6T+T1nf3PhEPYyM3ZvmGaUYXdc/39SQq5T/0KGl+LilAVQ2q
UxO1DXLzGDTN4q686UgefPvsjfKXQEl0XBqUwKzIacOBc9fdMWU5ztHSN01Vf6dyoznJYlHZWYNs
n7AyXPWdK1x9u+KdRkkvX3zGH61nu/gZllDKllJt3CiSBIwzDWO5Irul7v6ISM8Kulwrn/AWyweC
ie/U563Vr5n2RvKeIfOGrw7qgi4FJKeEJ8Hoj88gEKT1WlYyku9cmyvah0XOud0fPtNWB9zAHpNi
54LN/n0xk9zquVYnz5j+dGYJwPJmJnojustbcgkCpPpxY7RLsdHEPNFm4ZguHg0zxM9gGt1dDZIk
Ya63g3O+yC1P0vCl2P7H/tM/xRAUz8Pd/PWY+xodaT7xcAcvjCX+EgawRmpWIRafri9ZtdiFdH6c
aoTA2KEzbm+cWre94t68KBtcgmmHkiy/vVKte3aogQ+c8JKIFe0AColvzEU+jkFf8MFMnfVt73nK
7e2UXlfUbbQKse07r9r3EfWNpo20FO9l+kVvCHyXjeuBtYiQniGOwnStNCfGp3UA3jQ5dCcRUAz1
snxudNFGv+0h0hZ2NzDL5fNK/CfOPoqdx7wXmoVDxvTCRL555Ww+YGMjfcoYmByZx9egYqpW6N5v
4eLmUrE8Yvz57C44qpeFGz87zRlFBhqFcTJm4AaVC5uguLDodDRPSi0A2zP6JUbskyutvF5GqaLL
DhE17t6cyoVpniUNwg+vDBUdEP3HcU569Vw9gVrxVg9G3G4JgzyMoNI/U+IdsH75le2nrDFChyuZ
jNY6du59g6FawcKhFB+/tn03hIqw6yKEh9K6xJu+pjTtENhimNiXIeqiVAmaL0WWM3X7kX4jqc+o
dGHY4hOlC+M2gAqtOSnd05dmBbvEU/R3vC65ifGqH7oS1ciTlt8F5C0O+U7ylNmmVOihE3yT+Hce
hP088YGY3Clv7s5y60gxBG3bSNCkvJqsKFVtJ+aFegvlORhjVlZaCtzfrP6Draijk4Spyglp4jXk
hMxB2THK3iGRLaKPAm7QQtFPiKvwg9qjK1U3Uq1TjzueUR2X/rMPzMVRVqqSg3ysZozB91d0aLbf
RMd85Iv4a6m14mrCc2QCnkz5sf1YfYesSPBuGW2r/6AuyyOhfY/u/l/iF+PsHHgtrm6WwOLq74B1
xJIIvvWtola6iCn59lDgHMCvjbdeg6qrNHvfYUF5jC1p4zXT36DkNnDKhTgsexw5OyD6i43ABHyK
CJiKY6t/DX2OlALgU1aFyVn0DXNGFPi4NV8C3h6nxL4PXoWwBDb2v41yCAUFg41m9ds0xMwlq0Hk
kOd9lbuhpaHvvaGo3xItYEtOwIZH8lNEBhNehXGomDTzkUOHzsGzaoRLF1vWkzKew/HjQnPBaYFp
uqEroDpnguUjP918adrAWLj3ApyLT31TsexAnzJgZPxd6MdV2JMwASzloHB6kTinsPcKKQP2XW9s
ZaYwsYpefM4Zn688dWYwFN6FZugycccuXkCyQEW0h0sYeEXEYKZJg3OtZfsQFW0P5UOJMjGGDnoX
LO9898Lcx6CK74TdFludubqVdATQmo7ZNr63PSgMSGmiWn5WuxpFyr+YfmK7xhixULhU1XyM0cf8
iZw3hF8gM1uNm+Mog8A05BL3Dv16/rAwYEFeztiFGHEHM+LH9iRsTU9nge3/4kivdZV9YjS56zWd
BRHBz0xSWvUWFfIK0pI2IrCziEBfN5Ea4rNo2L1N1TEjsE1B+NDSU4jMPrTlpTIOI7o7XZtZk1db
MfYahxcbyPWWBrKU5eNk6P8opE7usF0inZkFe3g3I57gtgAqNJ7WeELSceXEfy4lSJlOSPptZgsu
2cOntpq8eZtD/sxpEmwh4/BzUJqoJf71ZIu6hyf5dMb2G6hrQcTNbflCrs6pr0HVQjCkq3KFIU5E
d9+2z8vel25+3UQlv1LNvuakQeY7VC8cS1GAEt4FpuGT0FHYeDdA6ArIfO39+AyZaXanOAgUcvCI
wNhaN9vXz5rsCStDaD4Zb+TOo946SjOvoEQcHXnrQahAjSznjAYcaR8HIk+a4RszwcvKfw+kW2mn
OwXRGYbWgR5fK97HbUPWH6V4a9KQT0V+BRoVIZKiyHcOsMDTXCYwh1vA16p733cG38rHSTYW9O/e
jn32uL3BjYWREc1IH/N9xSvvShy5qK2kJmvBrNt3Pd3JZcTmVHW1xYYX37RPTn6gKMUITfpFip8V
yWyPPS1kUIaZxvL599wjwZIauaqjCGLm5Nf0WNrx9KCFEhCYRaMCbZT5lqPZnJoPeDjsMTtQIWtD
dyNAZ8/xLYFk1bNh4FDBcx3s8nHPvuRKM3OQqdi5TksL8ake5k/+joL10w784DrwHw9DmQae0Asc
wuGwu852xuCsTYQcXCJ0Pp+SnCrgpM/cDFyKxo7tZBCJhop14AShADess4+j4HKHADMk0r8wqya/
LoUB7Lzrg+6mZmsxlasX/6bMgiLoNE27ku/Ae3Fb8mpO5VQlwM52JP/c6ZiFarLpRY4K+0f56Avs
Sb76+FJKluNJ+dafYUz9NbvjlEDZ2IG5SKN4qz+Mx4cYH9Zw7zjVaEJV6SeCk3giBYnIKt3JElO7
dvbpLTD6pcaxJEev4tIlVGLJ224NxGfywS3AFW5tgkBFybM7gj649T4QOaPQjVqdSz35SdFMPN8E
8dy9F5hJJtbxkChM84waI9xHCKn4Dz/cgFIq+o5pSxSoecygoYKyWVwqrP5ST1mILon2v4svx/J/
LcWLLMX96Ull1LxbEAOr0kxIFzMI0Y0vYTqBBClxzrsONful6Guq2/t1BguV87YYnj9KTnHvv14b
JAlCbDFbeqDVVhB2dHX6fxPx0nMz1oV2QFdw7BV0X21/lunOrFID+/eTw1sp6TBL7pqdUcNv7tTF
zWJIiQcBrW1IgDMBQ9h5Hg/cXC8B7OJh7cJLRT1opXNwYx/Qro0J8xQILTqZkkDLNUSB/LODMQnD
IcLaDybl90f/i5jiTQ4VO9g86sI03p4ZWer9uY4Im47Tz3ENL6rgOA4i0LinQRNGD575jBHs3Vwm
zgiM/KqzMpQvMtCpPBotgEI2BiV7Qkf/Nv65PwBAsFjHpFIlN3+2Ze78Rx0bIwshdIJcpQ+eTDNF
BxJglvT0q9tVnxUGZR/O+nf7OR/n4N1ip77Nw/6MatA+bYe5sWlY6rj8gv2ezUizlNaDm0syO0g+
DDrlM1jhBorV0ETzJuWcw96I2INRzzkd+xlaBqZYQFTMZSgjHArRJkb0TdqsR5YIO40yk1NufAz6
7JIrx/XjytY2PwR4H3mP0+zEQpUQ1qIuP1RRhfBlZnYIZw++dwX05g0eGaH6okh2SdXUbWJ9lt+Q
U5a/L8jIwsHmr2nSaHZWkZJUnH4bZASFiwsUOoxSDejPCLo6owwDjzjlDzPUxw3WCJj3kfM0VY/g
G9udup+GNZtofKwgRmNe2A9vFnIcoZ/fMPTAHZoa4XuZNK+3IyMfmQAERu/1i1HAqbffTJdFHMjI
1swyaWqHT9JX+Bgg5kl+whXf2O981rI/6o+ZGUjCHLW4d1cdwve95zt2OwYjtL2QVcwnYXOQWwbU
gecsiTwN2qrAJ5z3gWHvHAPeutjCV/PdoNNYtwfdSJAFLKaIO74Kx9WUYb0wgSMCBul4oOamS0xe
JyjvrCRc9eogTCNiE2RdSdMguQVKXk/vyh7b7KarigICH3SzB1rHNFRGXgICMEqxt9CdOV+TS/cu
Zo2AY4sL5ExQs/izzY7LhbX0XsQHr2FD52GV2JBmwG7oYF7QHAIyy3hwQ9pqv50WFeMzX+f4xkjK
tWibc4HrhHMVZmRLw9McIUlW/PBsXFrS/d95irsWtlA/J9f7fpf0EpqCh52DeqPTnDE6feRmUz1R
Ge4p2MIVFC8NAmkDqnz+3h+ys0VxKp6Ix1gs0mFZiApyC5ledmd4LWSh6L7feNmC2S1QbOYFYPqM
akbBtlBnmlH7dLkP/RnYBBgamP3iQUnZU1NYzIINzSND+KofL2ydKj++oTdD9/A4TKIQc6zs11t2
hz9ADX+EFZBmsMkm9VrMFaFmvuv+TctAJuMO+00U8qpwEPpdcrSke/KmTeKFiv77DWM6XpqHhMYc
R/Bv0Gj6AHlqI+Km9bhIuuit8yrGGC7Rng3P5NlqtDm6GcZisfRqg/NRs8mtFbjmt7DcbyVjPbq5
zAgbJaRYLBB6ySwOxZzDhR5Z/ludgYJhahNKnPkStBd4SPLY4ncZoPFVICC1XeYZg0OWz3oEmyoD
7IReeHv7nWeCjF/7tMrO8xzsH7/gFCPAC+G1dh8/uEg367eUZMHsPQuVGvq2JMU8M0hRGVwZUnEN
qnBVADrCIUKTm+1MOZcWt0e6XiJFVCPDjHG96mYbZeyOZMMKLNJ80zkLHZOdzV2b/xgSqx65VFmR
frs4MXy/8OVHtn2oijFLQSJcBRKdMpsw0+Rofw14jbBz6PQRqHq6vo3jOtBPTypvVf7j2okGtSvH
KYGq6rLRXg0h1MAWlHcrJ7IxpDn46I4q9RgKjOWxplESLzbLw2XmV11FgFIVLf21Tayai3pXQxXD
AOYujRU/zJHzkG/DVkm4vI2pvLSea+iWdT2lnBsBr5A3LpLx17eeEHPVFgrrSLVPNZAcLrmsxVtU
eRkBiuLbFMyrvNZEMBQe4nRXmQ+FjSevPnPTfTCMmFUVofjzWHVxhs+xBNr5kPUuuDDqFEkDxIp1
mFPw3E7wbfM6dxtUYrRGEvVv7CK8PTCNJSoN4jL+2HXKz4tJTPMcDeCFoDf/B7PsOrCPDQQECYnx
zHKBadLyqjZIO2JdKmOZlDcXuVMIw9NgU9qxMmLZUtURw0/80AOQZ0XIhqyOGr85detnM15X1LvC
YNtzzMLVJfkRCHQ5dwOrvXbDzTUhD3lWkbJBd6GvSEFxQg4fHH5hklRdsr0V2RVIrBU8M7+HRDbz
GrBGTIIGAsHsDl9t4tVktT0vvcmbr7XSEt1BI+YJcIkMdEN6WYuvFs9jq2H6nXJfKvDyelJYyihy
QcY/A1J5pAj+O2L9mBI+TNJ1jCqyZ8nuY8AS8jz+SiL2yvugI1JPBeG7xOko0g8o6Y6GRQwN7Fef
KHLAUg71fmdTX4ADyfWQRIeWlqmYQPcfvLqrVjx6SI3chAywxcPzKeNtKXijLSUB0z1LPr4e71YI
xdu4No9tQfsx68FD9YLCMrMl5frAWzZmzbjH09C2Nv9M2AAexbJWvAeEcnqGBt5Ywkgm4ir0sWyx
IPkxx+VJN0qRlk25pHi1eLnrXokvqbN+7wEY6eUpNj2tYswIkW5ws+7M83wohMocngSDoDgzKcMM
Iv3L1ao3d/l8lSeSd918fdqXn1BtxseVp7azFDGpOZYaWec39/r595B71n/zTJ348x+wjbz+cou9
ff5LFAb/3PWqI5sPe5th2+EIM3zFPA5Rjc8gI81LlAhjxLXSK1FpOEc7201m7oMJuhnG1tTyqx2m
I6cQPZOD7CQSwZ9XyjftItB7lB6WrxUNI0e6elYszolb/c3BNHmrupcv9M2HK5ib3tTIdAdu9Zvr
yY254Gs5mB5N37n1syEO66CzkhtDNj+jhfLsJGUxF+FMl5DoDeudJ6xqKrd22yDrNC8GHXAFEJ94
eihsW77e/ajsPaitivetcT6H6NC/TuP337a5g3RxTcRP+k8nzYCoMv3KhMb5RlxMa4KkMuVs871x
IUasiAaSHB45G17HNJOdLDPnE63y+xJl82lwCjLWwph3gnALdlUzKDMFekVMaeE8kuj9Lf0bhh5M
IOB7reb8xTMhtIvy6LlkZgQs47EKCAxKV1WbPEqIt9gwfuzwCpKbMh4HOjfG7DJ532QT5ay257ns
qBZOTHcoaS7aZGF85fnJctn0W+91oavUlqNeS2KhbP3G+1gRtsBLl+deu9URCf9n/ZZgJBu3+APa
2P+FUHYfSjAQFljKdoAuPli7lWLJ9i5rB8hghjbBPZ9Mfy4Y+BeRED1cfFS1F5yCCuNSHojbzaoy
ZAFFlb83/byneB1SAgkvqNLdnE4gcByCpIJze4zaE4bqbLMeTH35Pr5GHsqK7Jk1Vgrkg2LFj/4L
lerkXBLP0VPhPuwrZsxvhvRmnHRzhtIH0cSHkMWooSJ9IlxEc20dxmlbONbN/ykImJv/RSD4thl2
DHjsdxKODslFBRm9B68A+92OdbxzikJsv2aDbhM+MzI7wu42lgwa/3ahxrrvUaXKoXsx0e810rqM
j9UPeamPMG4glKOyZY84YFNmQ5NSAz0uRp2GDeBUiwyBTGC6Moh/AwNUn/nCwsNAOKPDLQPm/LOj
emD3QRnTCM5jQLymJPhCycxXNg1Gh0AIjlvaJ27zfhJCnZ8MxtdCLW9do9iXysMJsBfoTBgFZca0
bWyO0HPqkdCVLbvjgaKG9kNQ5L60OsZnn2QjtFOUZPOkGm9R0r2J6dGZ4lXDkU73uYSltS9fxLkD
ecTnY8AqFn7jHvWavUcgHpQ+83BPYI81QKwFtDVc374TylvHgVk+y2QYVCtIMjuMAnPXnVUs0BBM
3lrpE/+Ps2gymCVO18pLdp+69LlE6CyRTpZtHDOPNptv1I/w80lECnUF1g5U0EeqP3NRvBOcAwv2
uyoOGtdgY2VJd/MsWz3GZBrUqBJfoPRRFrUyvwQLOXKrCnEY/GmA/feBLXGaZ89CCFTDr5wtYFPU
RWoJtB2SHntjvGTdRIBr0/5M3rRxgjvRoG9yF+OtwG5ipHb0rCbCFiu720iU6YYW0LgzGBsJbvVs
b5srFKXCNGUC7rzbEzDgONSXGrZ0CT/mu/DAkfatcrfV9WmN1zEGJsuetSXx4f9RRbVuweqkH5BZ
e0sfe+dkGSMkZ+fKuwSpZTrS9ki9AA+Dbaxj6sjSzKmafYBnNBougo3vReMLIWzBH2rMWKRnGLat
RjRjxMS4v2VWNZaMpagQyFNr4mmqtfUAusXP+btWBwP074zVAKkFNldUReAHN3FL9Mu1oNhq9Pzl
VpsGr3+4Hw1uYCmkTpGOYzNi0whF8OZFhPa2GZ08xsS1WHQ/hj4h0MrTqFV9V38pTU4WHJV2EjhB
R1SLSEeK/zyHcw6wNDpSV4S3vbMei8t4pUr0UpPdg17aSHDvny199ZgUVbf/9rrT4dDnI+I5xiiZ
7ZE2Y3GFBrDiK9Rwx5yGXrrxTGYyRfP9mX88wycgt2O5otP6aULigMTWYbV7XSBtGjZculFy2FPw
nqHTMKL7awK2AGlfT4JueGkT8SnfHUQQFIZWlvRgsoq6dwbzy8iC4kFKOYcP97FTxC4IPJHxvrKQ
CGn7eKXVTP97kcVwrcGzIg8uG9z3Ml7g8ggzVrvKrikFwnBIYosnKdsid7QJwbzV4gOpDl5YcFEa
EO6CLjBBM0PwiKEuTmZyWCHQEBcpiyTXqSQ4l/0niVOPOL7C2ku3aFH0hshpYmPcORVhGScAGing
LycpJzjzErcBZhfXQRpLomvXz6BtLMpNtGqxK3+43c6VVOL2+uBgJ7x6+SHh/bBcaJW7Hkd/lBWg
kzIuJgG+qLzv8kt/NX0EK+tAMmmSEukbg41IWknkA4deVQzX2mvVInrxVcPyM+RM/QPbcr3erlYh
dcVSvN8QwHAIH7jtVtcr2Kan3VySSVFYYb4pKIfC04+Emroc9hkpOhvc0GyCFbRPbrC4Pqk8uFgV
N9SNSGDEG8su4y2vpbSFon1J+L7Jm8GSPjWuYjTFLW4UluRC9x2Ew2wXSamGoWdNukw2/+HFdTSj
wAkjB9VLqjbVwZYNpy5PIskHcIvN3FgeajnamOclTS8VPyg4o7QotsRlntF8CU+ks6ZzxP39ZOB4
AeWeaTnJa5gDyCrtCxCKIPUYqiIt5Mu0VIsNjEBsP6vQNhlLmG9dhz4ReGX9d/CXcrWMkeo4tq3t
K9oYfNcK1MfOgZ5LQsBAUp7L4l/rzwp7iObHM/I1tWjkZ1Q1NPUn4Dv8d4YxhDBt4hCf9T+8PXh9
m4YSIiVx6krtEqXJya5PiBqN2G4GVz3oBLJ+4EeDtYjeTfHTTJDC6JC09stybTKuOcEbp8DOQxuR
w8hpMSzhgmeCdqqlV5RpUmIgI/e/rSH58Y/duJ2J63xsygeyWIsBZ+60m8+9Ud7Kubro2UKFdKH0
F+Hhq/WzeM+c3jxPEEQWuvQ3PWaDy2Yuzvqw8rg0lnH7Zzn72Qe4cSuLyGpGLebs1lZIrqVbdB+D
czLvyxCHcK0p76uzPSlCmkAGxEiYVRBIIJirsSnMpu63qeGwolW8DJ+ttGweoYtHGLDLSAOjo34k
cgYnNfKgCNPzIzTq7503ltLds/9bc/U+pBmAirn/rbq6xn7MfP+3njwYNbjjdcmR+XGKzcAkBXuF
uooyMDxTCi5lH8ITWAnj7LFtJZZbmGxB6gVM4nXs3NWbRNU0X6NCBK6fyn+ZM7wJ+101LQzQCJkn
v7wd2EmiHUHLgKynWOGzHR2HHZLEHhgotPPW3uD9zhscHf8L6QquU466RX3aSIY843dqSxJM7AWk
VaXWljlMYBkbqwtwTxw34VOfekFdDwMdsrg1wIZKtrEORAC/xh+onwhgxFPwVd4Tis+iLMzE3a43
OuHnS22PLypA/otHk3EaUI9trAE6N2PJnOCb3aGODH8gG6lO/jQxfcNkKX8nTTvNVzAldE/SXy+v
Vx/8iiT1U+liZCx15x328i6n3tF45RTczlhmBnF8HZ9jBilcMcTlC6frwDdtqRnsNi2/CDoZ1W1E
U1ZHXk36bD7BEfhcW+1vxGrUFBYd+s/UeVvciueUtWMhPX2t5wI/RFJWu96KqcjIhrhrYC5UZK9E
sbxoPK4gCh56mSR1dWMQoVw4m7a8DhnVKhBTimCxzZHuE3eCy+bn9RSzv6fSMVn/c3aeDKjAu7aA
x0c2g0bGGbbFAtmvTIyg4UCOqnXh+NKAMGrViAd1L4yGFqvPzjLjLQK+YGzcZnSwKeidUQ383EOH
zV3XpFh+oerf+eQzA4bzDv66rcDheHHCq1QKP5F6AHdD72n0ydnOt2WquxcA19yLD2cw+19fnpXd
d1tm4wXBYJtLSt3lENw30h+PQab7HQ6vpF4LeFnlZkcIzFbCgkpM96VvS6uM6MPdAfERnkdtLjsc
Lrr5FDFtfHK8ImXPlraCqmrFDskJjrfO9xB8Vpgc3kW1isfR6Dq/qd+i8ezfGvYCRrC46NdnxPu0
2B1BtPjegoiv4yNjMk2n1JgNrJvVYAmieewNvMKzbg+kpei+3dtZRuKsdKoYQa4Hd4/J4E4Ssqqg
N4eQ1ySsIg9hneZQQRuqvZrx9hsXLJYxHO1wQIc8Z6UmsZqdECOjM5xW8bVJmsN1tXslpMFHHjd4
ywYOGwfGzgncgPl6QRnrFEdYVa1YgfU9PZmNY/17CuDX4QisXJG/m7VuYII/K+A+gtzJ2tDwEVnA
wHQAtUQPUDeFrWNbXt5rBo4S+ZtGdHoSqoM4s7plzJaM5CgX1na+i3QNjJNompplVoLR6wMk/JXk
ug1KJ4wmxrMJXOprW2cLLXnoh4ydcTCT344ksQmF1HtC+ZvJGDNUAkaHtjLVAXFVPoLDrs5GrNFB
YzUOpJ0M2NXvpMFyWCSg9y1l6G/g4lRDb/wR9mSz+I5FAgYp8O3cugN1eiofsC60Ddwse+BLl8tB
MDz32axck9tEVNBq02vXPM9J0XXH/khBrckiV86vWVuxk0TxEsJh0wcQFXbRmHii/FRP1yClXXWD
DjFyO7iOM3R3AWIOruU1eV0Vk34rSILunDW6fKGjEHXjXKL4tkAcRB6u9i1ELX8smsEmAZhKUiHk
h74OgWz1fpWJ40WSNaaYPoxImxVHGQ+dsxqTqQeE2kjNInPrFdwHF37tbrIyHSW8yAfTpHvqTfnP
eu5QgSgno0ydCyoNsmCERHZ+vTY22Nouh/nT4GplKYY8C0xCLmd0s24EXe/H35SIIEFlvI9Z9B5b
hOV+QJSQR9u6yDiHIW/ErJhu6+YOgOYXVgv6cnp47vNn1khJFCuQegucwFd2NlPtdDVu8VDWNorW
rFrPu1H8F+06Cb5fMXYnP8sfMutnpg/MRwsq2MIcUFCekJj3sXQAyWaMR6GEmE4kFm6xrF5qVXwA
bSFAWRg8wHKvNRustfmq8mP/CTWfj7F4x24/02B95M5kRYc1BgQ6oysm1kJxtaS5I2iP5bqXJFCb
hUbm8iTkSvQqVCVea1A2F8690i0+XOMnkKwegR50MJlrk5LBJBK3piHoTaHuT5gPBCLng/3NjiHR
fL69vAgyBi+YD7iscve6F+aTe97nef0uqaQJxkQT09eTRCxJxFicK4vDC/G31D1ZVmj4dI0vbSxT
9M3Bby2EQsX5OJJuymXzs9ciuIesMYl3bqgEGvjlRxkfT1y7d8BwVRKRaStY8kCFmjm2WL525wUp
/pbIkcEvAnAi80vgIG02adW3vaac3KM7ww3ybwV7ZjZjSPNbQdr2b5AJqTNlsKSZqY6M5XbIsb0X
faQpl1MWYJrb8P31w/Sa53rlTiJ34gfvWJuhV29KSWaHmXa2vbfV7PAJwEDnBTmHCTbaUfSsiGt1
fCY5vdwXy63fZpvZZSu1z224mJxnBlgKdYlPyDXW69dXPNA4NR/O6IEobjW+UmcXKZ2Q7+E/QjJ/
mbDQFL5RassTydXTw29dOXh62R2sHMqBzAv/tROib/VEVhbyzBs8aYVHLEMSuAv9mXMymXwZKZOV
cg1/zkKXwLx+YmnCS4gmrXNBQXUeuHQXtOjJpqu0JmlBcT23HKiiYHSgqSU1M6tJES9Nrqbpi4Hu
9iMxG5K12NWc/FjyZ6tRIDJvPlA/qKCF7NTXpW7M3mc+3rUcFvXbcQ5isnIYxCWaJG+gdbqGNhD5
HcdUHRGGmwnk76bDc8JRfzw47h4lxCIQTdXoXDgVplNTh2UGjxjSwyTxz34jD+MTyWSehNjlGQo6
HGzTf30ZIjhV4MY+7padOXK00poGoPo9uX0013B7cHh/9FaWIipXA6P914VzECZUchx5GHFSMW/u
N3yM9s69WuUNok2Rk0VplCFrQiVKK38k0ICaYbV3cPBclSWgZI/uBOASo6BnKh7LTgsyu6FL9+C7
M+uZ2RHBAELZ4HJjU4PoguF4WFtje8GMTuyRB/85MvK72/w3K3KmD3KlGQef3ZvsAL+RZEOMe9l0
dIDvwUwBMlkPcGw4afi5knB3eVNODvs5FYE+mJBfYH3SbGngMQvbQl/8RRrD/IYy62CW7LFwwS8P
PF7qFRlICWkRV/4ULAlQ90rD1sPWQTnAgTV5e604nc/hdt1bFAz5hjbpn1r23dgBPrk4Z8ZDvzRm
uYe3fBOQ63u3SbOWOsFXhRwfMCB+Vpbfyrw71J2mHAAspFqoZu9MWB/GUIdebH4u7C1h2MnqMzIO
rCa5FJvim65A23nfFfXC0DmpTaFKz4h1tEnDjJ1wUntl38gUwv192qwIr2KhwGJLklLGKEvJhJs4
Vgu5INmLx3VlgR+a9QhlBJqPhCz03pRpBlXqlJCvGAXFmLFfOjBpHltfqD8qUmNssKgDEKhvZOVD
Q54nZInCFyOW2RhqTKLDJ4jqWBFX0nB1sk2VuYfLECQMR4p6+VMHGvkMoHajaO0jBOvZ1x+Af+WG
WfhpdXQJYY3cxYezj3glg5iJCbgYvVl8mgxsTpTt8f2dqcXujUsYT6W3RT0JQkmS0s3q0HgBRBr7
JGEO1LeinyIiKLneU89u5IvEQNQwmDDweskfqsktEMe5TI/npuNidCPjvjZhLfXBdMYXwD2mwFLv
DEgSEOtc1mmdtlMdRB1tuend2OJGfrV5ZvsBM+nlxiMjTmor2Ha7bXOb2IzLfGoE5TPFrlopOrQW
QL2A5yRdJotxAYpSRU+Op7GVX6OAmJiOXoU8tXO6A6IUX/srU57Yp6CvJ9n7yzVdUnUAWSB6XH8u
fFNh8iDdvV00t7ehU9y5940ha+s1Kfi5FxQrOU6rBYPx+zRTyotkWUu2lpv94xhnEFynD4AYXkHw
4woCoZOl+aW0q+Yd5BEj3PXc2IM8HqV0Woi81FBZzhhCg4S+6/agzGSLjW1/I0aKYV/QRnMeyfmg
oHA2nydslAPqip5/MFjjQEaFTYtdhw2nM05Wg9goMCZcwBiGdB85/Bo8lmzZGuSHjmv5Y6f97J1T
sxetGTnKr4+yrs3n2rhLfW/YTGh88B56a8rk0zdBEaLt0f3VMokYA0e8VnUctYru6Sz5hFgNiYyZ
6knjmnm5G7/sC/RNuHg3x7KFk2ijvONK++TO7avm3+zp3PEVqzDYa/IlSGlb62IrdVsJVXgcY4mi
wcAxgD83feJg3bDwZNGjuWTID3kWNJxOKxAOcmZdPEcCgVji88cVmOrtEANq0aSG73unM1iP8HQT
C2qGcv6WP82Nv69qFUFtTCqwCFW+mM4JfVH2+vZeyWpYKr2Ew5lnTSj9cwk6sPXHymQn3sBevglC
ZC+xfObj/oes1F74JI2NQ6F4RAw3Ete4iFOvhdGDrmXsxPVVQZysxWQVBoQptgIqvuHjtbUmrCt/
MpG7wyhrpFn0S0L1SmioV3ibF/3Go3vM6Lpno82IIEtcJ3+is2VEUDSOqUGThaBmXPXuHndcH2s9
t26hEPDbIFkUOtp8W7CVSpDx0nHZk/MFkIviBTU91H8Pvnute9ONiRNvdMoj8+fdzuu71EHD9z5T
B2ZPV5kYrA+AJYxpumiD/tABFiWunP++trFAGTXpS9P4fJo8twlcdLsjFjfxK58JztZ/H4KPDURO
s9aHhGFdk/6Uzkn0EmOtYSmsNIuJyngk6sd6M233qNh7+sVjvJIwSygnuARnyLyoPRaD5lWQ7ijM
9hhITHso9PfJiWIrVZOz07XmcM5++21nWTGWXDtbhsXg5vUKITqIfZrT4jJkQJ7P9Jr/b8w7u9bc
tUlb5cyL2EWsT3g0CUupGUyJqZDrAPvfF59+0SHq97VRpZMEm1t/+OGzLnm40Ny1G4KPWqvxHOMC
S3elqnsJNVhK20qoy74VuO4r6tPog7eOz51FNI3a3A+sxhiFerBIHc7gOxAjAuJJXWm0n6N648Tl
OQZPRwPdA4IH7snYlQt/NjlgZ9w/uq8HlEGEAxIqdHdFWyrw1bGHuto5Wdq3tsbDvEaLNgwetCi8
+9uWF2uxPZy/e3EKAHhbSQ+/vMPDC4OF99H2QEnd3D3qTBrSmmbWqTpHnJTL3GeD1hClaOcEntCS
CeA0p+XIsnYjKcDNuvkkOn77mGWcG/sxzQRRQ3kSj38vlnfb+vVAygEu/rirLPPyGcelO7foLOy8
7ZShGfd5qP6jjq45FOfLayHBMM6Y8/XBVZxNVwl5nN2eTzWKACZisopKezsil3PP/08CbaVTM+S8
Ch4mvXsd0yfOGcKdeso3tlbG0FKkl3jSe93Sow6V+THglmfwKLYME+Xdd5B/dltBoUYaoemSlb8N
TeWv92+bQl0bKYzowh47oQF3q0CZQsQYomYMzgbs/xTOfsQRilm0XuAuSNjgu0gb8ZkMV/Tfp1YQ
zA9UzaugFe/xCuO5wUPtvXd9mJXPCYHBRlRoeP/dtvd8nwVFLrQZNCAQCQ9H0M0LAxAVPGg0AB03
JeLqLxHtCH3JdWc5Ugl+TaO6t3V6OclB7FJYYDD3vQ9igF9y/SGdnFkAknfN7zv4LQDZp9SspDhF
a54OPx1hfdIjBSzr8nVe5+xSBbdN6C38uEElaVQnuZnFvJJ5toNIxE6jrNJ5HILhU0XjShMmllch
I6R2nbkO6VcfWMhlpRPdWui9Dqj2qXxHtLCHmcsV58kC4rbU/Fo3Es1zwYHIey5LIOGp49YWoKju
9bM962CTWW1oV4hG2Y7PoXQUI0/GxUBPZ3VvEDgm8gaFbsWaEzX5DyuOLhzcWvhMeLhJ9VPf8HcZ
wiuT7g7MCnU3iJesDGMeTICePm1ErLNn/yUfwHkBDKLyh3wx+Z2vzkom1WhvAYyONl1W77+TVaMt
hqp6p4zgu/aReA0AkgutHudqdfj+l+ajVR6TQMTYwj8+f7aizqfXZ9n1WfjLxdyqJaKtbFCUHNOq
21+hyxmC6XSB3wvvtVmyzdJaSKRpxvnJ1VZaJ3lv0H4f7tt41CQiv58/5b8xTanIhmfvJkLVOxnd
wF7+gj1zMSC6lSIKqI/3oWcokN2Qznh/xVEx5FewDBNHI7nnaPPFwP9qF5erEJUtZhADPBE5+l7A
fTNi/ecR426NmRK//5qL2+ECFHWrCBpbS8DJpkHmULj9jemwSDENEEAX5Dv7PDiMtXQxUjGlH73i
tYskR38BVnxLK5D0qu/tbqWl6srRbqYyHpLGLFiQMLd6/u4HtQxWIX4hqo3tvrSmcDAZ5Fo34xeN
/NuYQGG22qBbHPhYDmdu7qATmbj91sbqkU0jIAVNN8/tVMuQdpiuUf4J7LcM7lXxqAm42A0jU61k
C3RAOfdywpgHid1h+ZSetAfIe/vhuoW53cDUFe619JMJd3NlrwCSt23Eseno+AN3iXrYLNKTp8pQ
lT0mmoLEAkL14Sg0J/IjC4RPmW/85Aok+nYI7hqbm8MHrvvbW1jhypQm2LwTneysdEPP0Yp3QJGP
pOYMRn2ZeKYDyEdJQQeB4SX4S+rNtPVhR8D+WTAYupHABXjPqNSUL/CdiNakbkLQLuLk0ylNjFH4
Vx5qd/i+NDiJ4+KimkTkwaeoHKGuTVyA5XEneRZvo4AUr6N5I26nAyfrDHVj1alGpkyhvajXqlkZ
4v7Yn32NAk71VEYAiyAaA5CxgyY3g60rjQAFh0wNPIMvi3bC0PhS5UGYYoHNJY3PWnqMukK/hrnp
Ux08LQ0cviIA0H9CzDuYC6Gh5ZDF0VtOuRosO3DPJfq7guRgEU1un6qqiKTPoZKBpdYuSThd5FlY
mBEOvPmZv0sL/bO+g++2mIUpcAvYMAmB8qBIS1lvftrxvYRpDsORYeWrLvx4zYw/irbGmREDQDvB
xPd6kiwQWTYSn9HMwfBQbaTbZjvs7x/EfMV67SpbmYfgHoflIKTqAc5nev/BbFqWiLG8ytR9qs6N
sanA8E8m+bG4lbzp7Y09xyV2P30i7xHmDkOEoPL+EG8bg9A50FP7ivGhUXLaSW/lUjO7Zo7Wyjdp
nig3J5ETDVxHmO3VADIHpc+/1weIOcYPYFmVztavWd3VO3iQGtuB+62K1gqWfBID7iwUoWqP2dTh
fAaj+nNG+G/XkSVLSLFars9FHjCWm0RJSJk9ANclW797EnDfvHzi/Bi0Bx+NrBIt0mkNatInwZSB
xACmzv8WAydvDl6AOoSni6F4kU2WU2L0AUIUMN8nU7/2ANQrFqUvCat3bVPcFbMNkT9wk5abR5bh
ZKP5MJxHWJOWUSKHoq58h9BsrcQojnIAVQ+0BrxksplRRSlPgoZuc8lias0o6DteO4T9YGnkkA7S
1GnKuJcvpoNvxK8czzag+/LIvUonhzes/QU+QnmZYSfm5KTB4D873GU0V4SqmgqF7rEwl+ef6Gu6
+Jri8AcL5tGfQ2J0mm8qw00KULrkkOFFA2rdARtE7Vt9FsQ/XAPWicr38AEM42Xvm2VQiASzXtdu
vUAoPQrb+1tr7Dvgt5jTcCdmYY1gjPs5eWiikUClsR1x2fliqMmnyZTf+PdevJ+lAB99S4FXFMFZ
gjYRfnxRFarV1izd410lVH18jOaExFeLB58psTY8Lv7daQbEverQDNFWbxGO3x01qMIjY+22yjqj
5xTH1gilYPnpyMisUjhTZkXsk/xFHKX+abzcpr5eARbkYUWK8/Xi49ofVQdAMhscx6Zos4cFoQKK
QcRtMFbJDo88gnQPceRFtyAaUYopye1mhi1gS490b4TzEXP+8yjbnKOz4ny2c5Ou4bbaaHa+kG84
gDn/V1DG4ISWwrjoG4lpqgSCUQTmNu1Aen2tNpeCWEn0j3IYnuKx9e7cCZNZ8pw3iCY8Wjm1/w7n
UPUvgD0QPJK6Afa9illAxz1g5spYxuttO5XybvV0HmCyxZ3k1eeG1fQG8ncfav/zIgsuvsUSANP2
CJtlWXCGe6+WH612jI7tP1DMApVKhGImmD1VSYZa1YOPQRfMhveW/BM5X4uFq/S8Ksx0xKliTdnA
RT03iTzn2HtcMD0+hB5YkTmLASkOVKtm8lBVL5dCPZWl+i7W+1BS3VbdXoLpmavS/UtSbhOO/hi/
UwglBu2gUlJhFsvg9RKRnmoxsfsLs1mh0RlE2mTJBlyqKellBNEKJ4PSrMywIskiA/6iWEsOm7na
nF2NKZm+lYxmLTdImPTIxu/G6LQ/txmEynEGSlnSNecDPeOGM4dEnaVL2J7UToNuq1UKRuPPG3Xy
aZ+9BsJZMT/4JdUMGFWAVWlOGH7EMWU9IvJ/D5wSmgA9qWpV7r12ITrXxegZsA1+sR84bAuPFU0S
Op6nk+JWBnDYiRm+OzsvNUf6ufirVBi7vj/9FYJkzkCLPbWsr8vc+Z1RWxnhq44VcKOU3HZW+Woz
t7PKuXiusIs3Z/PwkMawZQsj3eZIq0sNEZflcs75suvhU1/GcFFPqR2UyNnMeLPAL6Jrd/e20ag/
j8hIqna6w4G82m5OiaXcdLA30l4wz02F6RK5SH62qEfrEBOprDaH43esOVcWzD682Wjz9TVEKwxF
iJgpMlK9QdmcxsStSR3CY+Y9WQkMF54mALSq/nRUHggYEH6lPi15WpdqzIfwC+Y3Ei/yMO5NgaEu
77aYpmy0BNba4Ecr3cCn/XfoL6xp0NIIUlX039xn8rinFA1yHKBIN54jqZ4HAJXg00U8iAUk2TPW
reVdBeBmM1ahp1B6uILUeyb/XRMES+PK1elg0qhYKeW8XnYGZZZ8qwRq8K8NfR0aRIKZXEvBkFWN
jSTx9MaFYy3ypiiaA/RaI/M6pc7qIg0hC+XQG8i3QUY4bsStQK8qm604tEX430mmqOEwddRpNtTo
NELcLiPgYbBQ9JBnHQOz0/IpQRYNsux12bXmvm1X2j4nlDQeHNtXDg+eQUSXLV5z4vSJDe9677+y
vcSyA6DGMuF0nJVsQCnjgQk6lUCpvDcQfJUQhw/gWzJH2Yg+ia9wHfxoO12U0A2/ki+3zyx6h7aB
N1c1R7ohqWuOmerwLfykYG218OmlMVA9AFY0RWLgIFMNISdkRmHtHepKXGN1G7DFrIUI8MS5vFum
3xxjm53cfTdekbQigo2aCfMdpt59FnEgNET2YCewo5DuvCRKBzvrfwfVvuvsXDyp2HpFnNVr3nVg
815lMLwUrGbUMBKKeJlYX+812JzMZP4aW78v3oNDCYp70upRFRDYQ75hl8qG8PDs9SzzgpiSvQMC
JEnU92y1tRcOCGemI+t7WAfMlJXUpNwkTSw8Ezebk2lLHTWA6uQu7PJUKwoK4ExuBW0TIvidBOAQ
FX/fzFXLcj6uIiIWoIzdAbpSnvm+CHhIIGJ7K7cFBq3TjduIlZjwqXwpoHCbXPZigj17eNYc9T6G
A6ft2MkGxlZ8rUKHkBAE1E9xaGv55Gur+akx6iWpt0La4ebSh+ShBhO6eb0fXQd5imynuqvT0h/E
v8F5tp5nUe6/NnjyAEw8baTEjUFfgLhiH+DJPm33IhpfQoRNlZ/gRkm30Qzibgtp1DkuJs7I64ZX
/pWoJRCUq4Bi1V0tSjSaZc5CUvCBo34cLG3FoZpLhipVy/8wW4JP4qpDuvvswU9hSsee/VSSHlRe
040DApAP1Gj2bicb5plHSc34CdJFKBr5fMy+4wr4G5CWZTmPZ2dXo3L++jTwiWOHKs8b5LnzhSpc
AjSTqMbKpemF9ZI6SaQ6A5JXfHhRV5WQK8lehVWwYBg9Ezx2tAJTxPQPdQ1TT3/efvtIp/23xa1M
K+xZhE7VAceLQHI6BM52A4K+bEfsYW2INKd3oNIT7CVGYRwfLq+Xk932F6z6mFAA0FXteH82ji+v
IfdnZQoARzvK3XZlGUdLtcIytSySHvx5gqfjOVP52QgQHpUEGRclrk6AK3k9dlYqDy0W5vzFqAqx
Bbnc7DBGrrPLg0rKJbnHKGxaZ2U5aE5a6ohHrI6mQP5hVqlsim04mu3XAK70dqc06UrUGaiRHWJk
r4G16eDAErstqWT58fl4skhtmXFXn8GNYB/7jhdM31RYUz2RT30HO73VO6IRotV+9RrxRcUC8PPb
AfRVu0yIxRLvvOA0QaGbX8Me9dN4Wcj8NQWvdEhQB/MwboQ5kw5V1zPgixiPbqPcJbXV433mTquN
UxW80P6kt6vVhkVXw2ftbUiE5d3g/mdp6gnWOO3fBr3gg7ERvlaXOuTfQqicirzK8n4JhChNx0Si
3Gfbj/HpAA+xvd24q608U+Db+P9V6YFhKgSb6tvMsMPiESyP649t+9PKQg7h80EW15bRDMGnug0f
7unk56bOP5oh94WzwUehAKf85E1xkgnInCvNgTi5Qj4xnPOVyvzGSVAb0YHEDsiRowvq9BQ1i56B
mQyBz7o6n58z4NGYkzvyHZDT6kxoPtwxxHB2AaGxNz7l1k0NydTwhpcI5gogpWQO3KPdzHSNSDQy
J3FyGcDUV8Yst3utaLX7S9EKkJ3wCwGIZWU2LfUAcPKwTZhJs3iaW4SFJ/NI9a5kslGuX9zviCVz
Br9lUCsj+FxjJePBISHcV1FcRO1wXQvXIgooMqWfZBaUEdoFGVvoWkY8K9GLhzkPnpnjuZaYwQnv
/1z2qzLXTo8bLhEVPkmDre7wM5SljgcM7KQEHyh6sDvKal6ZPxZGeNufhD370SUfrqsKv7o9dZo1
T4Wqq6+giljUWXtyfPZ2pYe1JsNmZUgrWPYWeMSPsVP2USMwvpnRgwPFmELq4UV40dqAQ5gMG+hj
3tHaTJp7xIErlxJ92KJfiANdnhOg03tYVsh3zK8z5zsK+41oiv2Pn7/3uLoSUHnZnEGlAD9fMODt
zNFswAZRk/MFJvORCP5YcYYhULpnbaX2U++pcClwplpVZc9e1FV5kiXgQjIKvvdLLuYJJueGpvu9
yN7YPUJYqdNmeHTODy02zX/bMNJY8MrvcaJKHspM7K3XSV7wOERqQtvk4NGdbJFRh026a65VP73p
JIS1QDjNF/DUlynuoCRWT4jZPF6lSRfs7WNcFNblCUq89cFw1Vre4xEtmCQjCAgJJKMv4gLDYFhB
c5YxWyEDRC2UVUFbwl2zs3CiBJlOb0Ce3SF9PL9ds6My9OFyG+RisYIRbFyy9Se+Apung+yM7PpX
vD43Mjc8fVU2MBS7EyV1ZQCW6wTVFeWWd5EHMWZYIKYwd56SpWwne5u0PULJ3ByVhDfMfN9JlkLW
Y8ErTRKmPv9KlaE6DLlSJuULbXeNtzSmamkJQx3f4XMjpO9qZDhb545aUtAbz4TOnM/XWvWbkIXM
jx7o6Ghy16YeZleoATvPnlolN5OSg9ALIDMe6J5Eaq2LM38Rq8UZo9aClnXaMe1Z8QZuFKY3NY2X
rUXbv435qxuRJOORT7aR+7mu3tloOvw09Uijxm3/O1XXdOohvOe3VRtHsKc2qCLDnOBpYdJ6+Psr
jmj4Gx1yCQhUJRQhqRObsEZ7j04e0toUjCoyd4Zo9uFxFvBG2sLTEREjCIToxIn4fXnxy2E2/cvj
XZfV5eBsaMjAzklJPDAb5Lfq6yfRjEU3gJx9rv803Po3dpXcbvBFv3ksOv9lvijqTDFamdEqpupB
hS/s7fqFRjAIRe1xlTQ4Zuv2VC9lvJfVFzas13HsjoVqiCcR3D/zp3xXvvQGiYuNJ8VcQZBJafNB
l03Eo3SquBGWo6Fyhzp2KI8x2x2N46jiHKwAiteEs7hA0WxQ6fAOYv/BJMmxksBc5KXV1tOSpog3
YjAQQmFbWqa17SRb8QTdHqJ8ynZ8EThf/Grv7s02dVistaSHxgQ2axkiL44W+aBIDVeaYJDmWBOH
fpHl9TbXsCG42SAA7b1Hs5+k3FzqyjSlAer4/Ossm/lMpqMe3rA38L4m5/Dy6aedESNwcYJrhDt3
PJgR5sHdzopiRVgEEs7jg0EzOqrrgEiN3cEUB2P5NSc31dUWr1HTGl2F7TDSTS8ogztkdttIN9qs
FpL1nmIqtPUEEkZTIsdRJbIw05xjqcVWEgCtY3p/C1U+04k88WjihfiJOKk2Mbs4idLmd27BBAeB
jgCVqHyCfz3hKeGIeei9lYv8uWhQIbRf0g53wyJpa9L9RIuO8KcY1dIBTyaVVVUOOQEvmlNX9B6a
Ir/f1DetWFKr6aYMzDYQDrPbmUT4mTiea/9XgWNpMMQGUu28pCORmpu274dojhM77NUfj67ETjLq
UhFHbLp3sWqsZqhQMfVsTJYDGR/OVp9SzhvrcYy4Wd++60AV9s0bqDeNlV8P462HAr89YZNYsjik
BdijBxbuDj7iq5DkKY5X0Z/2bLonKuK+g9cuitza8D5OQfiZoeVMt/KtSdbrC8w76g+3m8q3goG1
Ap2ywLFHKpZEBlkSvbmzNooIumW+RQ/0R1Kjx8S073cXI3w7hfl3O0pLxkc8LQ8WL9kZTsVIXRH9
cArTCVDA1A62CdVHytbmJymUx76DG9RutHaEexrTdfejGZe7Seg0A5kXLgudbZmjE5hYien/pnIz
WfBwYTnz8lGkmW1kAYXf3HvU9naSdaVhf1AB9lfiZbWmPShTvVu0g8qvsdoUvQ7Cj7GAT+l3nN+6
TXQyfD+ROHPD9G3rpoyqa69604nLspJaHC+qwEm7EiJ2/+osVcDGxOSW/UN/GrICrCjRXPi6zH9K
o5rjQklokvamud+4Zzf6l4nrP6r6ACkdtAS2tE7SHEnSCOmfVxEyvppgxMJERlXjnCefG3rbUbwj
0oS+QTgbIeONCOulgpRoXgGsulzbHMkKycGF7b54GhzuyaWXpVJ7Xl6r2lXOdJ47QdwNuQlXrFjZ
5fULQgTK0RATL4jT6TVdkBy4t9smNqesRTR7dY8DXhuUwTlKZ8YXnsDcG36dlmQX8PtNTf8BeclZ
OrZnY1Cqdezokdbud/kj5vPDjnPsMAZzO4aH3q1v5S/GBS4I7rg5RW7rnAxB78jUtwa5X9SlEXgu
9Xvl5kV416qSQeqR4MhQsomcGTjkhyUAt8QJDk/9sGtlvvr0nXS4roqNfPGSwfaI02z2Y7pTDWOO
U3x1CdbmXkBwxcs6wH7l/EHh0V3IzK2MwiZbCaRfivv8x+ibC3Hz2WQJOnBnSqk04D9XcD7WtkFA
+MHryb5VqTwazLTk36ehcIlxr1FhBoIzTZTeZ4IHCJ34WqS3nW7gdlDOULWF1dNDfPIUbD6+klI1
lS6oDngcGdD66W1m+9TEJVl2HOi01trTvJKP49Bf/gqngio4HL7g7iys9d+YRWmKPYVWj2DMx6gI
tIywumiO9mloIIGfzXJNofxwp1uZidYxbukRxqypZLC1CiKqKJBItX7PeBVF0VCfN6JJ2HOGIC15
N7fYc8t6WQTPkcnDXSVKp37iZKFmM3SvCBXjcoQSzAQ0sd3GoIU8/QS+wVLJaPlGWv2VSyObuntj
nMEpJVyHiJS/LPMkV3j/py7CW+MRBEUUPDeNmXZ0jO8oc8XKywi8GvLPFkr1Nt5cbC5MTlEzrLxW
CKdD084JHljGSEI1iUx4vIYmHpkuXRfxNGn+QkV3Q0kKUB9YpHpwLajo7Q/1/d2pfryScE63XWqf
k7XDzooiNhA9yq89b0bbcWW1D044JvASDcmlWmgdxwJEEt7axQ+hmzbT6l9ubbAkWZp9zdIcED7q
OiCg7wjhqyZNOEe7EMCkTy6mVRKhVVE47lUt5L36RJBbb4JX+Ii5A7njAn2hfCrfSSHgyDGYRxiA
OF4xugIRCs2e1ZOITWM3fC9FM5UsuPM8P1p5SNdiZNPOZ1ncvHO3TLpY3THfMqdNWLLPdCRlHgt+
TdWVs5CjuWiLigrTGaPa59qvA8Eu9XnADOEhCktn858RUqLFB8n3XzEnI0SahRRKi5yVbiJ2+qpI
iULEmBf4n19Qdutn+N7QqeC6BHculKRnsWdMovswrYUW6vefYpQ+MDY+BOncMMTmjRl/NbIRs3Em
yYip1pn55Wco9nl3F9kDdKTqcy/+9fkbbI2wCcMR82G+zI8FdfdksxKUqCvQACwc3rbhXxg/iiEC
aOImGaKMyz0nGPgui7y6teEKcFI2lg+Y6DsD10NzZz0IVgESKza9qhl6HtPmGCVvxhnUNXif8uIS
p+mlYyx43bdEnU/pr/5h9xLUJZLW17MCI/6Qd3hDyJzSERKC9FA03WkBAs2EZhBo4yfEUweVTn2w
kaXE0DcG9rI0DJeB8ez7gDLXbiKPxe3mimoLI/Y2IwIf2txvlSJTkELwNXlPuzJjF8mlaiKFIH3G
C/fXeWukATV8Ij4d/i9t8/6YlZA7x6nUMyFnRHVWg9CDqq3gafBUg5vT85R3XUpRI09VLQq0gpTg
ll0b8jM3uVLFzbfvVzlLJvqc7WFAc7aNyfZ2j05SBKfhworhTajHmqZxBSkkUQwO5FlgIW7CEtm9
ViI6oWxeQvSIh2LZamLErwYZ/Fpx/SS4vpizQ+jpfCuZW17JPbM/+gRxGAdQOJdQdgrnIA9wODAA
O+u830c5OWE6eJBQMzqJ7/wiXgLsCsUCypkpFXr2D1dyzGB0vxYclMCxFte0RZ8haUHaxfL4nWp1
zE8ugJMyJD9/8IAERu4ayysyTGOnGISDki+xIXlxhIJdqz9xBsDkYJZoFjSkAUNsly6iH1LyLaxc
gOARniO5SVD/5J7x+YbMO26kr2jDM2Yh8dJO460B3kDeZfj9JCJsv5JT5SNb2JH2Cxfh1YV3474y
9QphBtuL+S5gN7d/CKfxmx5L13JI8db6L7S+CImBCUtb/2EP0uuoXt5fg4MNHMb3i/lIv4aWJiuE
2DNN7Q70R635OTegGsTNEi9/MKt1Y0UvIo9KRPnnwmswV9pLEKadBdXqLx5F8+zPhs4L8CGR/gVI
a9n2QPwFepu174Hwp1lbT56p3d2gB9+BC00qobKTHHkpFyky3HsVyKZ/t4glKVEqIRvPb27hQXLy
R4EDSUjnUVZrKut0MDEz0bWK3AI/AtATZ4O+oM+XxCxBwEZD3uammz6jZ2NUF2PU44vhx1WzLaSu
jy9siHOXQzhOm01SW9vBuW3awKZTk3MFejJyNJpva5m5n0/kKIIOg4LqUa1YAKU7YA0jJVXyYB2S
EMWS5+W+UJA6pKos9P/uV93i4/AAwcL5SVba0CniZ18YCCdWptoiSkmr10Pf2zG0+Da6by/a92X+
jKb+7GIx80zwqo7gocmZVtR9aVUpEocTMyzNMKKzYhKwkQET2dNzB1f9cnzZIy1zUDISNxiTj5lj
2tw9tjADY4LdzU4w/idSluj+t3ZL/9u0VndnUAwCacvgNCCyj7x8ysqo1ATzuCcMF2NOSkkY15JD
a505j/zwckIb4/3TOoj7kY58be+2WNBsOXdjHVRq/k5wRAY5UGf/4LhsSw94xhw1nhhBTdZphk2F
wA/AEdRCPDdr0QY5VU+bRgt79Blwly5KtvwdMn17PokvYDGHdy1g9l1mGBpdlDXacVvnzbzy2BUU
6AodLOnNf4Cs9Bh/r34ZB5aks0MOFUgbbL5Nwxiaibnh1di8Hbr5Wbf1a6aPzAX5xc4WvJTDwGTI
EcMs5he2VH4vAmkCtooa5Fof23wZtxuTUfl7l9IsWxDwpWI4/BvsA7qaInmcYaAvM8wQTGpEtKdB
qlxonFV6RaW0cAFKIJNssDooLbDtMIzDQQ1xSxR+DUj9/rCmAXrwt5G6tDcLql2pSFCfWqu90uSN
LF88ABjBiKRuFfjKfKwQF4YM+aU2HW7/Udl1x7cgXDtNaiP0H5V5X9Q1MFh3/mIUQeXxsRKRgvCC
BL3PKqL1VSZ+xW7xXV3Wnp+BEP6+iVaxU9V4DxZDXT9WfDAchpFoWvHU+L1sNGmJjyfRWZ2/aPEA
krFjjGv1/XLxkqhRk+rtQuukMuT9vxTfa69ZRiNvRnQ6S1c1WlZcqvh93QsWPn9Hrbz8sicubE8z
tMaATE1J8hWUtZFiEn7KsYoWkh3L1XFma9GL9k8FiPyU1QDEe52KyqZ6WKYNj+f7S/Y3XmIJDNoJ
oD0JUJdditmHpR2Ctw2dGZsDBC0tEDXfPHJbatGqC5qGDImzxzVrpe5EpZcXC43eLB9Z10JXI2fz
48MXsbP0XU8OVN6PXF3FPm9wI4mGdeLqbPehMD0nYRTgxJuxEKgCx5OvvSKk+9RDePnb1UfviE4s
QGec4nCGFUW12HF0ccywVn5s+fk3fHws46t8+qh6q8APpTCMN/T7sowbusOh9wB5QYMtnnYhiyEE
bvW0uplAbIhMT8oWRY20Rm3Qs4aTber49XTEC69YXvTUulCvRKh/jC4crbTZuq6aom9aR6utyNdh
bkFvjZXYkB8dkaUEIatxsqkVE0Z/ckB6vdKrpZSdNee5R/7F1vSnVq5r6nCZuWXjhW0GPTx5igSa
uy6ueliFR58xTNWAHNcY0gZvWRwXVlB2y0eGkvPRjalyc3+8cdJQGAIm4kJdP9IFPuTUOqDoM88s
KvMnWQ1cdBgNBScUSh71UxC5ZjE2yp6FZZnCrRTlUdUHSol2c/WmLMRlrg6auLwqIzag6UN5IeaC
jSjvn/N1q7GLqG+ckKC7QZoaQYs153DXgKYniX/rfapM/4y9DC/RPUv8NNzH9cytyH0vhQjuqfmp
D6UIuZjZxF6ScRS5lyD/6kiWDmbn0nDGkk6Ej6/qPdfcRkE3aKPO0g1EwmA+3rLeFLAMFHvz0e2f
FBOHz1zhNZVL8rOUK6vxzdUBbp8nsWiizkqTupZuPDw1WrqCHENIyN671REw6jRBS+gFEnkA+dgI
BJf/OfGiS1sExRYcrL0F5U8S165bNx6U7Kxo0Y606TD3a6lczhVrGF/95hXC6Qlpb0CMEFYfUNWG
+WpB6/baiFLxC3eYWl40jRJbKAeT1LywtRhw1Oiy2FTr0ya94X1opLq7xku5JsYfMQnDAfOF3rOd
b9MsILKFVLjdK6InETn0FfqkO/+GzsnGFL8eSkRGIz6fz28joUOnb6JqBx1MsZGf8vhmKzIyAdUA
HhK/H6mll5tLNLgLoenKJdpg3Pn2G44SOZ5nbnyq/UKcv/YYOytnYHI8eKfHQjzYaRxBCWPtk+lc
46t1Ov4AxWMseVzId3LfVVsId2i6J985NEmbu6uf4ViFJkd/i+GXiTDNMqchDfdJqRjTdyI9ZXer
oM1SVV2bP2nhvK2QE0L3hdthm9B/RanLUNKK7t5v+4eh6D0tcmc70DpiExsYbhN3P9I1pKosiFaT
Rc26usV4JNXfybIOpEr3kxDhC4oYruPf+wSDR8lN7Pl78xL0SgWfJJx6GhaZjUqxIVN4OrHGSIBO
YFoAMNY3fetq55wmwNuWwt3ypoHwsGHjZ2AtHgtibGoZeLdhd2v5GfV+l84N1MNU3+uKxzsQv7dC
zAGu77d77GLQX648DYtW8MAbHZhgGcWz5TIdHymQJR+6f3MwtesyGgYjZuJ8q/wU9ReA1i9LaJF6
nxiLa7k4aVIxWpuge5y6Hg6n9r1WMbyPbkJiiMGidlkcXduUImxkXQ6l7rdmohRrQt4j8vW03yYX
0mBz6p8YvbvIGtaOXG3T003/B9bn/ClQIwxmpWwYGXum4GzkAozv66KuV3GPTi5qhacQojoz1EqU
no5kU7bXeXXUJOdIFIS9eIaV3V98bDYXo4SM/2e2j+3KkY0xgNgjVEsFwJQ5tzgAFPgWjwanAPf4
CMsDnZQ5n4HaI8OLPrpEK4oJ/eEfW9TmL/PG8oO9+YNxgfQTwEaDDxQwU0Blyi/mCeiT4ZZsYcqo
0XYhM10njRzLLxhS+oLgoVDGsg127+U8uiC+jzFTK4P8uwAPmWLt++uRFUu3mU1kKYuMqWK1ehyp
VxwW0ZxmAY338TIttXLI41dFlZT9XRHuprGMv+y36ZDEHx1V33vATLw2XTgLhXDAWDEUy2j91WAu
YCWCZdN6PJExv4KzAaJhZgk0IVVds3CbzseWRKP7wZMF8Y+ZxTRPCteOsBPh6I+cMpcQI35CHjN9
jZh+x8djq5nDS3BkjUfQVVW6WUzu/T74SBMpO6lIud3YJlR02l7f171eS3S4EA4UtoIVpnPmzKFR
ShdOljCcyepvtRFQCaLSZLSWtDNvAv+Nxspv7AoW+vYPy/LhCn57OzgswHtSjcyLZnYSLV/Hso7J
HDX3v2T4heJ8lu4sdbnh4IqeYw57XVAudBBtLScWZLKpkWMutdq2zvR2Twm7wH9DuUa5gjV8amzM
rinNz7eN4VPfab6WTOGi25xSbk3xzMuWDKiWJrlcInRqOJ0+p6FJVy99cHZ0GQN+kay3mO2J/X8L
gmDp0cPeoYftmLPVDGhp1oWeMMuOu8oz3iwQKl7Ioq2ixJPTSz7iaz4uivaQaCA96AQTNHcaNE/g
SybZGhs4XeZCQnnjCPyymzprESYa7J+oDp7nJrq8m470SyCs9oB5YsC1Rvpc3C8Ho7gbdY53InTW
v0Gf9QUpy+3NGO7Ya+k3knEzG26YXyvin+8OJrKQtvVGRGMEob/2u6BFE4vgN/X6WvJTdj3B4eXf
8rVn3fofdbg6NpJNESnmkpBem8Fp4H5vWPqNUyEjv3PSe9atoXU/UHVA2w5WQM0I/DN/T4HyXTnq
74BIf+7Gac/ihVkrbPNMmAdzWnA9IYAYI8KCfXONh4qst6zYOARKMn4JGwkszHD3a0Ng1IOwO0PT
cSbHrDDTjoWAW91AeUk46caj8trafAog+2h27GaobfMGD1HfZ3F7h2+PMBmTQ1fI8eiD/jqdfUQw
Ij0GJbDdY4v6Hv9KffTcqMMSwKrLu/o/2TRu0HZuWIi5BIbEpBLGWsr5xJ2RL7sfnP2qT4cAZXkO
DwAAw9dUgf+ufxbJuh0hE4qM1Xlw0YKoKJbpMDnnkjB9wENr21Vm7AIS4JdTvWMmHLqs2b3qgLeq
A+Sz2pXAv82p5vwWfkH7CSMdn5dEncheAcqfvC7TdrcSHguKoj58xQbayaGFsKLIjFUoTWcar9Yz
VE1JEBxKmaRaBphqzpRGEPmT0H775SjgB9YH9EPDXauP850MhUWc0T0tLwWcNStTAOtb5epvlk1q
ovJU+PADs6LlqMOzqaPvnsBemv8nOyW6jXqJjoPAxuU4rzphZ7u703BlbjjDwHp+DM0/Ywn3SOkw
GEJiHbrVcexla++FfGZN7mBkDOAGoPbFaSdxzvSpNcqqGZIu9gmWwe4mHDRRG/dDNp8cJ/ZsIy6W
4g+tIoQvcnkFusigFNg32H36wxGQS0ND8+2/vHa5yp9nnP8isqlAuymxTuOVSG1V+eV4DMjwRUt4
J+2CU8kse2ImNYOHuHhD9IIs+2y6mf6CKQJXHaSQeTx2RJSZsdpoJjd2btTrCgzaEfRw7tRYKOXA
ejU/9KOP8gYL8q1zzY7Kln4uxHDt1ROU7f3/ESAiMld9Cyg36qjQMEbTeHrPz4p5dg1Lk0C3HxW0
jxfkI5z+ouRTQCxP0J8F+HB8BJdTVKV95L413H4sNC/6dbFx7VT39A9JhIR423ALc+TQupodyItV
9t9cHloawYveP+GaCILY4c71zUDXxIfmG/8NLb5rL54VZrD77gE5uE1Mdnkc3o+4bTIfICoBz/Wc
LNujFW/YTBecOoC3Ca/EGFlUeKP+EwDI5wRIdTrqE+UzkfR4EApUhSjQsPtXTHUUXkwixXCZq+Z+
bvKdqfYoFbXnCP0VliNKkHoYPTyuJ6X7kN+ynw+m2Y7mt/ulxurQEs5TBbB48X/pDwjlilA4fVSI
WongDulj4p6ODVJ1l/5MrsSuU15xcKqU7FyHIZElWTK31R1OlT8RCvWshTliSiyNTPFjSecmSBdY
zSD6BxemiOX1vefRIfnO0Kfok1M6lLy2i/LAJlQGvXxtf4qsTrdr0+Gn1+SBQHV8cJ3P0ZNcAcvU
99O+EPOlooD5F+swAR8IA8+VU1+KlGs2vjcSPQwe5N56jXMNO5y27xtTE27T/bu1kKshTGm+799U
NG4moNCLJhH24pB4Mgdhgwcx1y0oBosQm+ryYfZ+rToSZrOHBZbZ/J+I8gd03t9Bxupk9YpoHzzg
kxVXXfXnIG8ERvVql5ZsfG6AaaJkDwnjR3+ZdMff3MbmM1WSyb7ud7Y3pNektYanw7QJmMdkpA9I
fOXu6DT156jLo0xZ1eWzPSWzqUR5Ka4SwaS5ulzwY5xBM7VZuWtZDP75v3Pt4H2r/quJD6YETJtp
YJkua3IJ2FWQmB6GHACwoPjEaSKS8Zbx5yDu6+UjiflslhRfij7roIo/8QV6BMtbtczSxZ6hQE6Z
6+Tdw2eafzm2M6wdwUmtxwvQYBZERHGJPwohNtreC0cXLwiPrHTJeXe8YgvIes1QY+6jDDMSPn6B
qAHYy3g/neTl85sc5KLCritbx6cd4O+zzEDRla/XNq2nVO9Fx6NCYlWwRoURDZfLbxDEZwjOoo/d
/apxGOd91yKWecrDiB0+jfjkzRLRs91lI0GBTbcSaquUiRUdEHuMqipKiac5JEzVaabqYCT7smVj
f1a1OuQvJGcOdz3S5NHtGF5y/pXnHdpO2qJj0h0prkI4sXeerxGEr3dMqmzWYKeLbirh+aoTKN+/
r1jVe/WvOsNw+8se7IE/wgrGCtliSp3Igu+ofwtNgx1REfWgQahryFxu/3bh65ci/12pORD31pS4
RaVl9o+QUVgxlYQ1onlBpyJ3QcZ6GBCRozQNVioFOj3GpDmEpJvexuYJp/NO/oKDPxMNCfpw5i+O
ew9O6ghDBWCuZOCCpIywOSC01SNe05YsHPIoMnyhuhZLmgTJqo5ZDX0jRWo421DdhBGtUXUfo66P
U7MsNFyvGuLt4rJw90xB9jicWFvMcy2meS3TutVW8IJSn5AYHoQSAtwYi1w0yFQSeA3guQLKPa1L
a4EU4iXdCenRaeCAWP/976uJovtmZ2LY+837QGGl/G7XrJZ9FDZfd67EZk1GDekwJgG1Cj4GyyNy
i/q+gq3K3Jw2iRYX6T4K5E0gFlOB9TAhs5m7S/R1FcHJ9QsEbpxTh4exLDMt+HJzqyfARruDBl8o
WpY3Y6q6LNLCcL6xReeRnBi81KH11W/HfGHsJM1YvlEP2sEzcVNY4lQMBM+PHZghbMcVE5GvoBjt
HLW6U6e0A5wBnO7sigwpuCc0gFe/H/bIADwTE/nqdKwuUbUNJ6EAL780Ai8xSkPcE+A5dJzsrw3Q
s1kB4A4UTMRCPkbBPr6igXIKFZsoFXUHuDfeKefiiZoDifZFjgYh2h+ZgjLu3r7wBL1piFqvcF28
MPRKtASfVExVPgTvsX7/vzgnzfPuDqEO958xZxpJoON1qHpFxFTIyj8BukE83ObHFV5Ddyc4iVdm
OOsHJtO9YhVkDB86vgUOEuT+yULlfBCOc/6Buli5plsdFRZWBy7Luc5xuM+jBNPeXelR01NowRvz
yHE2u3JOYp2lnseiL7gAK6Nh9s5E1TQPpgZU3DHruW2OOZxHjEuQl7fsII8+KZGqib0ueTYoDTFa
XHjjsE6dMbPl3fiN2k2ZHguQI7+ombqQENT31KRu5Res8mUzJXF1BFcQWYWcS4xTuWwu4xsrnUSV
FIgXP8YFnihAY9dGZHuXhvfwUzEntDtq1VpUybW5piOHdoExWQQVUU5iygnvjd6sUu2cXvuueLcU
UrqqCUC+wpEx8RwJYWSyXXdlE1tbfCwWEJ2Jp6kOGxwyoTggH7CqdHrpVT7yapOJHJ8myTgkjxv7
j5KgD0463lFsGP6t2OAF5JD7XGEsHe0SsG0LyG/xelrKguR1edRZw6N2IOCMDM3k43YhiJaiHZxY
hBXJOaqVuJ+3CReUz9ibcuxEE/nVkhAcKLBPpQEmv0jFFZwGag+mmnwEqoUvyVGY8v6Cq0hvLsK3
r8LeYZwL9cXsgIt8l4O4kGSSkwzySxnsZjb3r/I40S6ENuixYk7CyFVMWrqmwxqIO+punJsPVIRr
A6EuoDO9KQJkWztA4wIvOfP+gBrNsCpp9Mn7nS67DzkWg//4GFPyF1mm1A271Fjmn15XyNFG35SQ
PLP3285UKDxHehOVlibREy7+Kc+ClXCBaaAm5Y9tHtpAKa0yPbkytkJt9sONl/QUX+Oehm2ze8G5
wh8Q3C/AqfdolQbph2tyX3yFJjR0QoGLv5256l41AbbqlAKHeyTor5oR/mLPbO9pPtAl23NOnJ/p
ji4ZIEbz8DYA/cr8bVkIKSbhrI2MNkIqa8RWKzdfqMOJmnfo4OLO92+JlWiUPGPHvDeeCAz2ioIb
NwbPqAaZyPprJvoxGvbUa3XGDs7RpJbD88pFozBpUG9QgiTnxH/Lk+rttQm7h1LzLn18pnihtadp
HZsC0SsfQBH5kgV8QcjO7xHB9sd7r4+dbDs6SNCtJZrxtdJF75SJklUmzKTwGY0ceGnfffEnjCjm
ygH8ES6YgOmdBFSQml7Kj/wJEIjYUGdLKT3Ezl7l59cUfkMsZ10DEnxzLvzVU2KtpU3uRb+oGcMs
tGPUHcq5wNqsZ7gNvHJ+9Wm0moEGw7nd+4HVKoZoDsIDwd5wwb83AOzWWGT9upPO+1eN5ciCFiXe
HrUvvkpENvhkDgMR8L4/ZJIn60Zqop0lk5RHIx9WoB7rwwl+n2iSYf3WEQzuIlqtgSsrFzkhfpoa
YgsGRUS29S3j0GEOXJP5d1QXiZ4tfbHUjR8Ve2Ffnmqkyx+pY0qxyPP2MwIxNuNEyBeUUSKS8bl8
5okZpAkZ7wxt2hXx1bZQ1SmJwe2p7WxfsD9xwSf/1S9NrVctXs1/IZkYsrU2aseptu2PdAgNSmF7
FWodlnhU//MIRtOPTWd1a9HwhydPhMoMLiKvVSxbYe1dglbrLnJlc98HnK7PPzASPvXO/U4B/Ygn
UOPRhuARzzKr2dxL/5KppYDq1ULGgGma/03hceEgDLsh3kySVchVYeFGQB76QEXTa6xY1uXvALvT
nm+wewwIS0+hGOIQhwgJgXI308Z4Vm+QAaI2EUgkYeINaCicT66R0VYnZSvaJuX0ZAVGh90kl5Cb
LJEQJ0yjFq5tjftxKsJseUgd98e2AUTMydzcuOrADieGXu7e478+SEN+5BDycD9LydANZcYrRu6q
IRZ5tw7s9W78tTeBH6RuhQVjtYGlT62Kh+HhcyBT0fsk3KDTbayrHCfEgda4M+phNsNSB2P6Ncji
gF/Okyg5M2JHK2ZFbAAVaBcfkXqBOwiCXr7aNwPlrVgP5W9n0IO61luJvgOL0jHNPOavfxaC29Oa
/WxXkNSGWkFjBuaqGj6V4zSr177JYP2CA2JrM1ZuBJeA7/+ZM8n0Vh7enztbOQche6WK+IxTnxoT
aWgU+9f5wARo2LrxUrZwaUnACKyJUJvz/JZSYl0Wm005TMMHAdJcMc+s93FrbAdBjP0VxPno6YCo
AiW0rFG/02EBcEOBQXCufyrzJzGbLVmwKe61PNO5VO3sYabWpvBoO/7bFqWFPeEOR1CfxJbJ6ihC
cZwXdfAQuo2FK+ZIuV+/gKHsSBAoBmEeSUSmciw9JINJU2+GY+mgXmsZgnHJpDFvNw+PWsgXovOr
S8Iy6APrQiS7Dg7K3/Gq0rmw5Tg2v6TLIsoFrYHs1+4cKpKf2nPPZDNToxfrBEyriMTKNzaVuuuP
UOLMCLAO08urTCuOyZjn7J1T9eSZ3HVXMjl/R+GHZ/2pb+5NKvAfDdC1b31NHGYq/PutER82LIzu
+OezCzn9Qhy4qdEfqEC/J/iW9qEU19QaSdxnnq0OJSGpkHm6QfDcmzf8t2bHLNtp49kqJxZ/TZEq
4+dI85/pCucWyoIEsGwK5vdQ6oaBLmDL9AEicxJFlWjMCE3xnO3XtFqMz+/k61cGoOtS6kfD+wKv
Exs4h2bD0kXvv/7NgoOLpNMZKrRWaJrCllcAW1masUm4eiwCmi9EXObZWABLF0GKnINz7hCcWBeT
UBJbSpXYcYM0T5nrA41zIkc6lcsCx0HV40tnu2JIlq1OHq7yId8Yum4ARtc5SLlLAX6A0F0IDruk
s+BcRY1oAqrDWgxbQWWnevXYTBjYOro1YO2BdIdgn9Juyfh/onciRyT9FIlC04r63/mgR1E8k27T
TVDALOTps+wGSM7+719zK7d/kzgpnYh/xUfZJLq8DR6xE3E2kabXieAXC8oH6ddm76iwpFZxwawb
C+rqsg59VeIGuBkMWhB8m8/vtZdhRDw/NQMUDPkqi3Ood1LHh0a+Lukne29it2JcJr2Z3nNQks4n
V7mUOtBUnIdmsLFijzxxSuJT+F27XCifgrQoUnBLATnZ04uzrAODdsKJfuWb3V9or4LTjm4FgzAT
87PrWO0ENHM6uzb4ByYHmtnhEM7/Qc5jJrBptO79KfUMoGYUwbmiqXRAHfrz81+3QSCaNDOCFx9L
ptd2TsWAucTeKZRuS8XPzyHKxz3YpOF1UMZ1TwTUxsuMkJHir5FIoX1W3PbtYvt2zlyNKDNp80vb
dz8o2k63rVYD14xTMaqHP+a59dFUH8bVF9ZK4+kHs4owDWk4uEA6anPnktTHOVEKm7OvZpX9pt+K
193uodmu+eX30CGfgnIE+fOlrnf0lT4rw7wxpNuHm9oUtRulTQEqTHLt3kaNy63CN7IOrrX62c0L
XIR3A+zg3ey7NDkWEH4nL7RM8dJ1VX7mY+wnvsIWXAW3c66wuxU96LNvw778aGCDvD51r7fdDVV9
aCDAvXbe+Ba6SIUlm003QCDWd59klUY0I7dI5RdeSlQ5yJ4ztbPpRf/8grv2Xuyhb9yWTj7M7uNT
tVl7hNppElJsuyhm0tyZWOw1l+GZ3g83FV6V2r69j1HNqC7YGtmvSo87jOOedDyKotapa5lCbkZ4
kWZ54A4SRb7Ol2lNcrq7Nj7CjyRhU05pEFBtHAZuXcL11j2HfiFaxGF8NefS7vnZoL5rLPDHOMUK
hrgM6QNNxThgNnWAEH8r+ggX8v25ApYzfJc272Z4NmczvkcD++QFSLfeY+5S8pd7gRP4ALLD8nPd
GI/lxCxo0KDfZb02GomqyatHS2wJYd8T9qHfCPPE5Hyd7liBEwtkXOVQ/HOEDw7UpmMP61EpIFy0
euEz/f/ETWe5/t/4p3tyQhWoz7NtgFH0yVMzUWPR4MSXaHpR6sPEj4T/BMNnXELpszYZIwH8d3ES
PUGamZJufO6X7aD8UZ4cZWDeGPrt/cCwDd+ZV8xBkZCpgGrSmjAK78O5KtnLc0e9/3Py7beamHqd
l+tp78R5+BOLoh/1K31B6FzPACAhnSPAtneEAXKRpht5K+OyCBWS/gzWRz7b6EIygGKi0HUH3B4M
GzHuqfnnWcpCL3+H1ZCL9NSsDd1BuIgCQ/x/5jLqpp2t2GFqe4a/csVcphW1GTtGYcHT1JA/rLod
QJDsZK4vP5oTnuB1TVDE22pNS+R8EZm54Mne4zVRMdJLA2kUiL+OsSipyaeoE6FJDTl1pmSWn/v2
OvhlNQj2WUa63myJU88yJ1lAe3q3pLKFEEOeMc8ygCZ5ziHiiMAjKInW64OFTqErNrhOlL2NqXGG
4lvR2KPMFfJpMun54qeRNluC0kyebRXp7Am/WRLW9Be9zUewgNBclI5zmznVoUmQ5c8Mwph+3Qs9
CHzl0vyOummFn9hTaxExNcb7EhlEB5SUzh+CTpwMVtPJyuEA93BHBAhNAjcUuz8MibbyRbsWrE1+
4B41fyuXjguJl8X+JOK8XLNJH2XQeOAqj/TuY3mUh8ap2E08nh9kAOVqtahAgjkJqdY4JdRy4/pe
Z2ZLt46Re6yS2ZNvM8rZCLSCa3Rf763kqqTE60h2VhAsQUFdPu3GfjqEJhHPCLSdnh7TE/Bn9Laq
H/sUhCzyjXYlUGB3+jrmbV5UMqXrlx5/nJbU61YAJufFsavpp16WZmx5Tt0SDxrITxY94UHByqlb
EgeEaQBLWInZTXwjUl8q4umPD9Z1EERYGp1644TwjeytYxttbX3s2zwknbQ4UGHPN1sfsy61662Y
XL7QhrSFMgXd5RRXHYWK4b22O1KnrsCBFzNp4BM3PERWJ7yXuckMEc3mwcrvPK2UGtMPQeU9O+HZ
b/MSTVr37d9sNRVfyBjXh0onfE4d4G72f++hbCxOq1e6gtC2u6lYFsWVKaS7wrkH3MKiomFKTq/u
XTHpf0YdYdrNa87A+24o+tjnLERf+B8s7Y49a4reiqVS/9cSVw16SrUsV6i83kNXB6AJFE6WS0jk
gPL7Xf1IUigHw8k0k6BSQBuoRqKBGUxQwWajttYoRc0sPV+3VYROTpyWlknmYRT+ihxTQC4p+KNi
CJd1XdTP0GgaNaCltlKJZEI+ZemvQBjAVdsGYTtEqQAoi4ri4jZx7HGtLEbVuAXYDfuYJku8/tHm
EuH/g4epCS7jnUrh3hTpAZjUMwYjjT57tguy8+hjnPnWL0a/F/Uk5KK8KfwuPKIv1gcANXe31Gxv
w0vafuZYmjBEFgvcztMdv8rx8Z6vsE0mqxJFZ1Gi5R8KnRsbJHdf994oWwgZdIxOHtdfXcCryVHH
pQ9FjiMJRVRZfDjx2RBK1JAi7tFNibCFBS636lWJ8dtOcxKp21bCM66lhdB3jx9/2ERAwzIiFIVv
bN4eWoVOgQf9uoZHTtDp6fzBkO21bWjriv+9uZVQxjyFz6ts5yZPwQjZ35weyqGkW+T/i/V45Cvs
MhAYxc/3ynPP10MwLysxc1gtezFKAV2k/f+l/Rlh+6XLMB+WMAMIDvEYKvRyj/B7PoXvw+EqOZ5l
qQ+p+gBm8DKCViE2lKVtrgolJxc7TYb2pkTZwuxYbSMkWwOB3/feNWEjBBVKUhNIgneHcKhAfLpg
Jr71n+4hf/Tft/cwu6LumFzhQhef35kvPXDCjWdwgNSoY3NZBGitU0IbQbbXaIl8BrQE2Nw3UELY
S8ve2G5T0mtTGSBfISYLCLz3tWnzw9cmzrTlK8crS71eqX1fZ3dcVRi6ZMfCWBLcnCpAaULWdnBf
OS4XB6bcppQASXM94ssxfDun4p7URFH4wyQwg05/4fyBcZdnUA31nDBdHday0kWc7qUrW95KN2bU
USDmANFW+99EmRmJpVd63cFoB8eporsqYPYrVUz0btpsV0m5IOgYpI8L1GJ3H0p/vubfUdXQmIri
s6fIUW+tsJTVLITPDh/8BQA8NwJ1zUMR4448w6Ctze+erq0Nb6lks0k1lkBDvjns9DIt8H7h+QbL
KolUeyqAqUyZBGIsxQzTpnLi6KQj+A0inYo2pC6sDHNP42k1gfvFdrTdi3hFwMqU/ICTLo9A7FD/
EkV5CB/e1mAHPE3r2ocql7hdwnUkjb3dQktyoT8iz/2uoMyfJxkAmCfnWYtDXYk1PrXNdq7DsqL6
nMfnU91DLfu01LkOLCl2AO8KSsIiCjx15luSBRvHc6HiHE6P3Cq1CpmjFJo2Av4j9eBi56gSPoyW
dzFBOoMqNfMxSOvSn6hA0y1WTBi+g3vZFWk5lqeRGBd8I5l9+vGyhANi/wru6uRhPBoi+9StnzZj
krG2dt1j+KfHRARImNyVneRHzt4MJs6W1/+ADRs+suSA+jei3ObZY5Ae5tGrrWPFV7hqPZvEPGnD
71m+3Cfg8+54H/Si5R2IenWAKlI49r9ml00ZBYrJ1gQLHoz3LWSFT08t8qKK9EelZp+xQ20QhEXp
TRctocwPG7/xdG6fomDVFBS6xXt2NP9nWeqwXtssNl6322WZ0z1MbJZKQC5DTvkhntqeCZ0grZ7J
3v/9lkdAGrC6ODxcQ+mH5Y7dQ9V3RJrm7nZ2VkEMjpagkjBlP7FzBQgHX5/kqmR5PXhKppx5qjcV
t7MFmCd9wBKcWPc3xoKWk1VvzfScKtCYLn3eeEseoceUNu7W7QUuNXcHOos55xjMIqmSt4SF7FbB
rza8oqwEnHyF4jjazzBPeJd5nTk18iYvyRSQnKTyfDSmLfd8RRBIx9rrH/ThiH1uOTfmeUzyh7E9
bxocyY/lu9tSkKNP1SajdbaUEhQR7phHbeW2emAUbjKGXUtZuP5bugxZoPinIzKcWKFh71d4ztAG
zSbDnR1St/4xPO7DBSfQqTQ34TGDtDqkMHMkI5QHFzipWv0x2vGfVdrmg0vfSsWZUF2+xMYiJ5+F
aMXYOclSJMf6NJE4MoUL9ecpsnYKA6VXCRPYtdZMBwa2vYyj9KaWItD3qO5zszvUv2PAXfPxt7w8
OXNneHPmmHXevDSf0YcwPozjTkokyE0PoxEQh3l/fymrRPU4rKAZeU6f1nFBFs5FOXUiOIFJeQ/h
c156AAZXUdqqa61eOgUc3Lu2ywhCH7owgIyYJ7PLiV2k/1zoj9EfKOGuJYnSkNzKld2fPCcXx14t
9vgz028bEZCzJApSjqSqiZSOp71Yx9BFGfZE740hlYI+7msbY6cWLagsv9eB4CMheNlluAcVNJ0M
Kt0U2rsPZvS+AdlE7uLZhUWdS0cGN+dcLdq77LaH/WRulEd3YqdJruMPAIvqP4qDrJvSGYOfqaJO
XQnlSnPdjLDJkohT97bTcXxhtH4KBN9sC5ZXWzw5r4i60KJQveKMDN4TueASzTacWZGcspg9CkIV
C1aGsk2BjX19AuLnwgEC17hefdrGGfHpHNRpov5x3xggCm4OVr7VKzcW9D2utk5Gk+d7PmaWzwP7
6lMUWLdiS16os0zisp91088nWQv1HfKEGPnXaV7ZBoAT//XxODxGsQqe0gVuNJBqk4gvAVuoEcby
0xmLvA0aUSK3nlqFnIbcAHJ1bj4J8naw1yYxxgZpJK4rWm/RCMPOJNbLq2IST8Whf/gVxTlqrkc4
Atn9b2Pp0oGNjwjHnabbos/H1tRFDgIP0E0zpLAj9EsIAf74Wls5AwjjZZ7xXrDX56C43qjDnGZE
WDQfxUezFT8131JWrl4kMQE4UeWNYU831PZwJ94czJ7u8HaNlIpbtmvqSHhFm3bvGMQe6a26OL94
FRO/BEGENWqRqBi+uwa5kThHU+FkoksklS9tVrxUq62bUoy7vsCUSb1hynzAp3GqQGjGPQgS63Ya
2woGYMOCaxGaztCl4zNHeweQI9VoExjyFxiHxFU/l4y4wfwlGESkUizamjhIO5rD2g0s2Zo+wJm9
hIC89MScyj5C/AqO2KevcPUrUTihv/hTRVnQXIH6B6oknFDbWQJt1+gEEgz+agPv7Ht5lBlZbILR
vyYfgVEyMhQoowCxpQAT5BrXogwQVMCSkpjPT2yuMirTpMlJVXdwwJfL1Zg9barf8XLgfLXwpvEy
326wb8F4hrNN5TVeqLWKdZD78SlCsR0fiN5wjOtryKezA1J7KvYyb2uTeXk9HAhpDMc112/4FCk0
Dzlpquf+iIwnfiWEDuopENMGMifRJljI1q09uRg0vi5PQI05AqpKr8j51MVIzb023R47p7OVS3Rj
xsE3Rnt/TMzGAuXmTY74WI+I49hDLskwSOOpDRKS+K1QzDoavv3ygic/d9cbwnmUUG/fR8NkUlP1
e1gm4jOuUOxofxkGKrQR9q5ZVJiKxxEIMRCtR3C4RJKWsWBV1sqh3726LoR/L+AHWjoC7GRnBlLo
Kzm12BcGvF5MIMW0SEXWs0kFsP/Fmh/2e5GKY7yYXQRQYhU1FQYstbGuEXO/pBA9dcJy4LszUnnv
+dHWATrp9ObbM1PNZ/0W31CU8gpLd0LFHv7MP0rdXIjVzw4+OmrLvugMyWPEv/Dn3H3colwNV2OH
KVOnbu4R0UEMso0vSh8jYl1fr6f1xZ9WiCkD5P2+w9Stn6yEiD4pyDVWgQsboE545DQud2lnXkMn
kE2iqkhXGF+LX++9sZy0aVgRV3ZQ8Yp8vUNBKF2jqGMa3BpASpKbaOXnppn/TSxiFSmdKg9ryiUY
VaSSYVC14bMXj8w4uONt5y15qwxGjKVdpSEc5IFLXP+ebMNdKnj/S3x8A32efqhgXNJ6+4yH3GMJ
PpodzPVpmeUtj2BDPc9f8tjXQuPDN0QuKNCRRUfPQsGlWkwnmSOEUUXzAn9xR7kN6G+Aj2OXBNV3
AH0pJdanayKlM7BE9AQXj0eQd75dBy4VNROYYWepTJ0wg3qUDc2qfSUJJXmtTfD+4B1MJ44X2KNy
Tf0ZeHemddVcQlD5HlfYTxxobu0pbzOXx2BmSRsYvVVE+59jyNMnSl99EFr3uwlaOePO9UEidyRl
LwPvDlAOV4Mo2CcaimxdRN4XtDYgrTz3Px0dGILphD8oRW+/k8xZKxuz7wRawmF9AAtYPQGyikTP
fbw3DjM6CwtPmcyshgjxAj6XsjbGYDrEFM7FwKMSDu475sMeLgo7EgeCKr8bo5bKLudpl6OdIRec
hYjTtzJsBsUtx6PbSQYpYk1UIuqChTvEmr6o9WAa0tbwBTSMigAZa711PffRU267BwJK3G2kLvXa
kmw69szlCL0j7FktWAk6HbcgI7bnScvsKhkeds97sKvU+fnuGZ6AlWfDMrYPAkH3cFXxLv7kIEwx
Ssyzex8asKwMj2zKNT80aClF2QcFa0FyjRPQWW+/pyzKX+k65CyKxxgKxNGVPJZuNjqDs1+k3hED
EiqJJ15ICXYeO//WE7ogGPCFrkUs6EgHyMMI5JPXoj4qvIAKdWkuGkLJmyCo/MGbRRlvsKjZl/Ep
pjFrmPrlAzZDJJQTmnNgQcptbHAInsS6g7rNg/UztcdInzUlWBp0P83kRBkp8eZQcJq0OFVyqAwb
t8JJPN47QTy8Fo+PdVn2G3dPigYbZMvMrdgVDRsR9m9XuQyxT8ofQP9TVGRacb/t4LQTHt14Jl8k
EYUIRGkOfp9nklZkjAG5oMl6zDuVm2Y8rD4aojHfROKTnwXdHd3MMMQyxUL9kx+rQnoejdymtlRl
O/+FBuL52AELes358VdNOFiCtlPO5T53zUuS/9z2nzn7V267I0oo6uivp3vFjERDdRi58wD+yiZ1
fCRnLdAgevSKTQts+b2k7qcD1VLPr6oPReVfRtR/Vdnx44pskFe6Ez+7zHaWjxwl3ZgdIy5J1W3i
67yqlwcRR5u8nxZxj2xtUmZWywv34i1NWdHmEMA1YjzGObsDFTDEeGHBM2xl7RO8uBzTxdmZ45Dq
ICoLmNv6TMrAZ+W4bOW7Ju6bXwBjbQvY73EDX+dpfhr0scX0Vql3rlwuA8hVrIgGSyHZ3fJNEw1T
5ZQF3GBk/NiYPSiC3VO1RKuPDdEVNwnl3UGoJ397MyrWzgzWzhZNGKsHNEx7cF4AffexyZus6QhG
KeL4q7YSFpvQZNwtcrOfsdafIsOXALgFhF7wtehpRKbOksYjNVzqAqWPNWam6MiVK0kOPaMkOVfP
cH6yjE24CBAnO5jJbaUd/40J3a3V7tD2FnRW4sXrn5sS4ifoPdTgy0csW4eS7O4yZDLrCpATTJnu
bqJpNglBA/odcs6PRBbWyfchCD4ztk+/IBnclnH3g2ZiJEXmpw1bMMkMLFnC7gLKopXVA1R3KHdl
FkOAUJabeb0pzRldMYdKCCWl+TYz98XFGba8iALT6uuVjQflU6opJFb7JrUl3P1ZzcRCMDe4oyX9
Lhph3Cnvuvw1IjJ5MRj81Qg9VfOMs/y2TYi5XWf14S+oSXulKwJb/cfRXev0RYlG7KRe1i2rrggE
ey2n7zqM9KVk3inoRUBky1NRBYzPK5x1mM2SJt/53pvkcGwNN3cgE4DWmCj31/KOgXmV9i9aIE33
ZU9ba3oooY+2lDEIICJr975ljCPFrYHiCoAp+awHXr0GJXrel4p1Ax6wO8FSNSovDqGDM4IS89ZF
2T0Ii65+LtoKZ7jD3x5fhczfDVvHULVGt5QaUgU3JJuZZAr4CJH/r33HTx4UeFPxCkCcGXYK4LdU
VJpr4hgjI6Aw1MoEACwRdtZS0jLERAemOs6y8aZT9QigutsEf3sL8ZaBJ4PIO6a5sRv36ACLLj78
uGO6GlND3BmmWwJxE1ibghSv+ua/sURO5pE0xXjuc9L5SbgAW4+qqZ4w7PNlE9cGXbgkal3zbRCt
p5FvWqldxxebuuO6lsd1b/0ONnE2ayAiB81eDLadVR/dY+qG3JJE0P25lNe9V+qjf3RzpiZn9IFc
wjNsG1Kazmh0aUcaBDo4/2oiS/CmCJ8EApymv0/1B3GWnGnI2i/0IHSlnRHeUEIlx3TdmVryummi
VB0zZ2+hPnV7bxIM0kFfxLk5oUvFgAVw+CBO/x/LGo2IKjmwDQ9+q3Zq4Xe61w634UV02IKDnYlH
d+xQOaWpcxodvd4RWveF2WdttI8XuOgTP/11BLBV3fo4Olx4r/5KziTxW8P1ur8iEe/Ia8xZynHN
bjZ9Nu9skloj9Fvz0F0gkD0rTmIOTXikjVtm5p3E3J54SCTRSbMxN19Oxv6+dTIrzmoNIUEjQmtx
HX1CF1iHwDdVgMVhIK1b8aZk/h7n2yg6/O+nlQuCoTrzOzLW9nf24GcBGV98cryaYqdi3uR1TRod
Z5nL2zZdQqzhu3Wht7lxy5bFk5Wb47h7AzJ/TMkWfkq5qPBI9ShU8IQ1nlei3VcveEwMFjiv1lwx
rHRzksjyOuiNBGRda+kk+KuYoyS6ETl21AEHGjU9W9xDM7ZAvquuza42DJ7YJzO8wdwV/WU/pPpp
fMvXzHDShnlt8Rv9OZJFmmAoz/ovQRftCGouQLByEBk7tc5HtnJ+Al9TkisVgOFuILJYJv/Merpa
ludymNqNxkejNdYi+bA0CnrelXczgxGtE7hqLigA69hpClq4eDlGatblzqUjgPVzHLAOxlW5JChO
7xrgJX++QB6dNN8pc46zdlJYOR24pjmO6zoIeghd21vRg4KGVETZ3lmohIMvX3zva1Es2dU41hGM
/JtsdUt+N7sfwDZ0SuFgLgCKFBslBdxi8YrRpGnHP3+UQlzPA/9s35NWq0RxNRDqTwHBOCercn7V
bsauvVTFn8nt8SX2hg/YZOCGSlZk1wefyLjj72DZKIxHRIrPPuFkN7N7UJM1rBWLjuhp8xC0NbDU
Z/owHE5RgA4A53TCuOKoGXN6yICVB7jPdKLEMCmTiM2HygINtSlwGk7s+7Mgn2YGGOo5v2/7GbTm
c/5XDKEnRpehYNw84sn8FE9xe6OveIw7E4Z0HzoL2yGhPlkkaG+89zgh9pps78xYD9ZqOizDS5RY
Ho7p4c3ivyxIjQ1k063b0Yclu7NwMY32hvdoHAT754NvcbM/wUenRUBqbRtewHdbKhdrpuxMpIDY
gsa2aoN9jmJQoyBc8+6yVJ5NtupKpgCdJ2MPc7xtAOokpncsRo86NnD0xRTRmMl6RYeNwNSW+F3M
w8bIE4gds/K688OH6qjth7PRGG/EYHCeYupkkUyP/vPvqTKqh1QzbHWN3Q58F+o7AyOeiZhei9cB
8+GA0paKYjR84uUsbKuFPxMEbenf4zNc47M5MkV/rEZPgPfD0SxHu0L/O01Q60I8Synue1By7XGl
Tj5aMdphTgEKwwQOj3dY3n+ryD+56pC75tu6o8yC/y3jtTHozlFRgzWrVk36+zjTCrjToHWsUQn7
w8v9Q3VehLtC9pvCCHCptMydJa4+GOHBFBOnqvTx90qiTAr9TNlkbXVE61qKGFciUyyS1C+GfugP
Sl1uG5x2D8R8pwJ22DyUyLCj0cxJsP131O/ouB7Ks4A81g1ukW6EzvMgL2C/FpqKB78EWqqG6c1j
AJns9ucvhXzbcr/mhuRc8iBlmyAzu3zn9/l+zIkvO8q0tSp11thoZCiIWe6yVU7pxtOpEPHziJyO
BNQJv9VTQ9B6hQK3vFUDCwb8buHJkL5nisX9A9lo8dOtGIoSpWrTxY3HlfxJi6tkosesKKXHE35v
ZR/Fd2ws5/IoZX+vsQPMTbqVy3dcWG41FEMQOOjslgOEOrtZM1S8zlUpjfuynpeS7KedShFNwQ7/
XsL3Y8ssyYE6jETXHcdjbmOS42C4dOTAy6ifDWKByCC6w2sCWdN8XGcm2gVezFVV/MBQsz7/mX2g
oPRJQFjJn2ErBIPWoHw+4iyysVaK7rdpQ4p+C22M6dEUrBCTBwAXvaPVBPoUdZ1HcaUMpmXcXpWi
Ebehha68X82kcQ0wDtT55sig6yArPSjkDIcoq7IJCNjWmrb9loRNZjnb4LaBCStsGOn0r34SUv9M
IHFyqHKqhbc+thiPuliOSmOEOP39G2H7dSL2o5Cfe+NIaTfsw26wTHl56s3S+2WH00H/ZfxKQXH+
CMOETuPmMGQfFfiFcosUT6ExmcuBiSMU5PYAfjodVZkYEClhgQSzsmRGyJSZRjstq3iElOh6PJFD
/sNps7NaPLHCBCDVM1Grraxt39daVB9YlaUmUmoK5tWLYYdPtgoiyUArjcBu9FdAdDJ3BSkhc+4e
RyAqJNntnZPupMJs2ty3Zxsn9tOfwacamRBlci2/1nPn0ocxJMrLOGN/LNdp7ynuNEV9zujzUrZx
j5lwuVC5+rf/hlwGLEkThVVQaHh02jy9Zi/PkbSk5vsNrDfDIixNYieMXEYQddVJL+0LB6szsWCI
SX+gUyTLYEKmebmE5pcA2ZtKzfPA2uuaifPhvq0Klqpl0lFBwHH7+dMFO+tnEfadMXm/Eyvnu5SF
CLzes9VUrWha/w0Nq+DFRX9STZUxUoVVvOFqeOxGhMC+TBfBlp1jxN+wtFRzZQM2XFdmwk9O+mtD
tXpz155awtQ3rH9Z9ME+BjG1iqW2QjI9j0ZFULuzfi7SY37xv3gW2qBt0WY/bQIFiU2ClHcAaZhQ
Bwr5PO24gYcXIvw0RwL1mD6HmTUmve3Lp6FZpZqjYT6aW1lFLbXxMR1+LHcii28NDySsKj8MiQdO
OZ2R8ochmgzZQiS5gD3qGbQiqpkBGZtu0WTLIzOh6oqDTFyJQvFWAdFNcHubi1j84Byw1+HHz4Xy
MpYW5WXgqBZ1ze9336P6QOcma3FdJaLOd+11CWM+rH0mR8t+2l82ZqIGnwXsaBr/ShjI49Oo06Qw
Ako+WIobMH4GiFg3t87sJqzouR/AaSn3cROo7Uto9y2z3C+MmOLwv1tVmpEEs3d4J3/Cyq71/+EP
JK+MovxA5Fn24Uohp0XYqd0btSa0tZLNPOS7Wk1zM2Q1fAiyPEWuetup1YKJ7DNlXk0BzzYFciEv
rGUTXVeyu9JSHEgSqZ82xNkW+GZD0knyQNaxMJWAXnxFRPT2w58vcr8rvnwvJcRxj/bbD1n3o+RO
1oFi7kRUEji86CgZsxHD1Bu5DK50X4zLqcP7Ffi6meObu1z75C+VAMAf3yCH54yKbOcGvcY0UgnL
GakCeI3NMnEccb4tof9msA6N+xcsJspVQneWZKhMVoUOKSrCygUsTl6w8IrFGtxLIny3HmIjoJ9H
Q63lr98F2buXY0boA819tZ4jfQD6jy4I48/q9pTF7YFsWT7YqYs09uFrwin799PAAjWhPDOftTZk
o50KyBfe5mqd382SkUdg2hjStSpP/BQLUAJp4dPccDyg5Zv6Vb0nQbDoag4tITkqYRfd4lqM36Ab
eEmFQsB98DENgFyGPIRZJMnGuwwdwanS1HQd2qRSnNQ32I5/JgJIgodMsPpAkm8fw5SDGsNIpQ//
jskR3N/4AhviKZ6XIHZ9OKQdSDDBw4typYzQLwKrRo4+cW8OOW/tn1DzzH2vVUbcAwHHvkhbHs1k
xsjdUZhkHiWmXtoQqu4zMJj5pmq6gl7yc+KezR8ool/7PI6xkg/rAI72WcsmEvq4SZ5i18VXiA0N
VlVW6QcoRvYRyxE9htEkvVRxUEEU9DyI8gYHaDAY3SGfQG24WPmFEqOpXXuL1Uj0I8iJ9mlT2IRc
IibCUkMGQN33puUmZWKbAmAPdloG5l/nQEP+7+dY5mk2CJkVxhKjw6BQZC711PeEX4h/d9kzCXPC
4bfpUriOuaFWDQh4+6CQWoZNBNbnrtgCAF7pBRAFkbUkkI5un6IuSlhBn5XJsU9bkEIUaYp9veoj
KqWi1/HGhkdPMcthHsgW3J+pR5HN8ZC3RcQGBVa4i7FHaRmYnzUtHHOGVyHv2W2n5Z/DO+V7IKMO
LDHIMx35gZo7jZYpF28wycD2IRRvItKpIfNmLXStpqsoBWsVlS8L1IyPuljfZttWp/lX2EACpZ5v
+qLRIMKoFsIGcMGXbXhTx6XXSNqykY1iFPkNLqCoNLOHEf3U18fCEC9Tdlt5det2b8FWnPS3sgb5
q57ChYhnOVzbynbL/a3rPXbjQHB7BNodk+Taq9ftb/5xdh/Ao8hJ/bobaK41wfRfjsRVSzxJnEcn
KJv0+wvOApVUu0Fn/2aB+xO7ruRLvW9PnG4Cfjin6VL8TIWptXXhiCvglKCTdTcBYEnYAC7+s90M
GFgF928GjhTkntxYbaoZ3X8aVgYO9l4XF5z4+Vy8GoKkwVNImJ5DoXjrE6qjhlIchnkyLp5Zb5d9
ltApjBspfjdBfrW2R/TwwER+s6ZHMN7rBMvJ/DtnWhS+uJTTAbQa37JJcPAIKz8mfDIE11kZKrmS
0qIZFV+ip8wZQXjYz1MUShDWUFU443Lh54UUyCOQNVgjMuV8Zh54e03b095CxkgJdYeLhONcuMCf
3nZlUyLHqWNXhVpnuUo+yuJQmIXyyU8DADfboA5QWmNR1Rrv93m8G9jKFP3sd6saAHhjV1u4egK0
ASgjkmK2MAM7k6NPpgqp4Zo/ojmzWC4lA0j2JBG0MkpNQ0227PpMd4wLIQVF1zLMS0jRlqZEQgNG
FRGdMLx8I/5AU/WFvUjN1+Y5p4T/BXUX7KkNGYqbyD5J57pVLIB/2OoRkGzNf+9vcZ/kZRvQGNVL
5v5Ltn/gXYPzAM2myW3oRaiJ3oKDwSm8n7kRwjTDH+DRJakzZcS7UM76R8j7Jc9sjyZmFUPK7l8T
8PkmncpczQqgT/CJNvP93nGRcvaAbOVe4huv7O9RDtInB2/v9trYaPk3ncmBa1/m6Ks1JMOzeaLo
VQR5bnnXelbyioiAx68XV2vE6r/KxSZSF4PuuDfqX+J3rIDVMXzFGqJUXJ76pmIX6gimUdfVt5kq
oLUE1wymRGOiNuUZvY7PTDIG9RzfVmF766QMOiLLfJw+NRMy01MSxhkCP3u1T7lWBLCky/PMnb+J
MEcGqtMpA6pDba3BQ+D2Oa9f/DLRoNWVfqFyZ6Mce1UG+3iaLV1X5kr33eRX/gRAXSa8QikLoiWz
Qs61T3JP5bNKcIQ5rvg4CtvtDSwLgNHRrT9CttwiSs6dcrJihPy9Ny0I0V4i1sGMK+UiQqtPByg5
AEMuVkSrf/ub+VllY7YDhuK+y0Y5/JSJUsznDjNM1xZeLFXI62K5Yz23jWmbJvWZJK016w+A34Mk
NRar/kcj8IHzQ4jXgtltptv931/15BKVbpCNzF7F/mlbKeRA0Qnu5eoYen23BDpbUgu38wbiCe+5
LcTqZTgEns8dbDM2nR0vvL3+gYmrPwAbg52twx3MKo/1DITYpPQo4Fqxbpr+BCpZlGfXLxskDFM1
yeX6/h65tPyBOs3tQ3UmU4YbWN/qS+DFcXShYELvYZjZOZPeMr9q2B3AqGx5F8Z8a5p8NHdTWp2Z
GccIuXm2BpjSjF4nP05bJPfJdDxZheNoZVL+RIREuEdZz3SfiALYsvZnmhigXoxMa/RataKrOm3R
yDJyyTvv5ilNsOru1aC8uhIk04wcDwO4ynKAQraB6U9bwVvdXGs/8Ke+sW94g0TVDw6cpsFFliB1
Q4pTF4VDCKyQ67bSdyyloCfXZQz650ACEJgKbATXrSMUZzg9SUEwjfunyfc1IPS6x2pkuoqk3CSW
Ro3l1KWM+1BHkOIPad+LAEwseIBSKltttj7lqQ21ydR/us35KD5tHmU9PXIUbSD0UhHWnPOcaC8K
AZ0qO2LYWYdtqR9Zf7b8i6lPaiYJ6pFtwTyI3kEH+/bxbWxO5vc+eQNp5bzAMNtt/iYJbZOoM7Mr
rh5s6beej9gPqssNdohe0yTPQ66vE0/rmvQzW5uot2arbeoP+kaha553JtikCMoAJJP2f9GyUMqw
l2CZ5axupjL0nb5QmUgLOxfA4dzYHRrQ2tYQlVjXuQSUyFSLd92ViaFaMzuER8liyhWqp5DX1qxz
P29ANWuNBrZ5+UwAUqSC2z8OxYwMIQyc59Bf2+hMMlB4VnkhIEVciOnaepy8KB+OXG3TqA3X2mCq
GnTGyzodKEB+3A0pd86OZEEvLmLtrgf2vO3uJUxPO6YzsPTE1Rq/vCGq1UUBtxifumzVJSPxtH0K
8qmkRvqRHB9vfkucEMHkTI5OXVGtdUR9EJBRliS4CKNihNhCA4sv+E5ObfG0RVWSEnnbsqRMlFET
PL1VQj22MZntROXsepuitnN5/cD++Lafp19v/g+wjGrV2bHJsNjAqJ8S0vgD0OhpPTbjorRNx2yu
N/AIdGGVh0UloCIRWw8Ht2wRYetf+xPWsP/hY7iUZ5t1uReSbeXGfox4V/lg2k1WYIu2wz0DqcPb
NVEIe6EqjMoMQn52BD0u7k0cWMzq8130gcewgYuGY9JGr1YnLzrIepIHcTkmdk+FL9sDezlEpbeu
ovumN55GGtkKRjJRLDvzGiJMgAUZGupG3OApHJb2qLAONbqOF/93QDFS7QYk4f2y5yCZabx9ZLj5
oXNeu3TWThzWZu3n1M8xpfpD5+/eV+Grxae6+ITrJAS4z+vAgrA+usv0TP0dhT2G7kejbr981IUu
ISLkWAqt66GpFdBBQPSeQYm+NsUEVYLgzZxaqrw55vBRXTmhDIx1feyLhqE3lfI2yQZpXGuQMsgo
ydB8VtLU1dPV6ch/aNr+/ULaGE9sUNT03cQJ7ePuIwvbP4c9w0rE9UuzBa2WJ3uPckqpQtEeIYi8
HaBXh9qqLqvuAJDqw/Yviic5bv46OhASTiFavBINW5fseHmbeX/9CotUpehiqZOwb9MmcxRsxpW2
Xav7KM03TtLo61mb/J2/MlrU0nIAtO16FKQXGu49g7yirrJrAeStEQ9lyd7xEA0mJKdZSmYLxxr4
hSn6gd7lvNtDF2i/eGwih4HhPrrHyatkt+TIA5qiyd5I6Hl7C1uSwJ0+F6lGBnNL3cEMF4zIjgtP
Tt3+l/TgZDvbHy/uKUlvzdMMt+0q9Hr4Afkd6klNYsG5c54y97/h7w8hiABKGKGK5T7EbfXARvtJ
R4gAwwB1M/IetR2wB5yd21SlS4Mk6L9bBOF8SIgzxDSrwULt1FMwEJggKgWHvK21nrNLNzhGuOPj
TMOQq+qjKz+D7bIzB5l7B7fuUsx33GOxfanGqpA+eaQd0hDK60yKTZICb+GYh7QZmqLGa00SEnSw
QTcVgesvl40VxAVvxw0U98wDxdBr1jEeFZItberH76nZZezDmVsY2/+Z4HI9APSgoWmYzhGtaRhj
h+3P7ibCJeWlLbzsv6uubBBBWwvYWOJODegy2ML/IYKJdhwHU6h/L+dAIB+DFyDLVujhXOedjRE/
0ePAKOewEb19AJOcKodmolSKQWTzEKzJE1uPLeDp7G+GeOasOptMLTi78sTBaM2Rp7mDu7PxflWK
bH3eXclf96OdfkyhKiPXgLRQlvFgTbTS1U+FgCEqmGHJzNJzk8JryI1mxXqON0wHaC+9xiqtHHe9
766sbOBHkoH945RPz/QtfhigxrZ0BHcAVNM4qGNcgpnUPScHAZViuPC66kb8XyHCTwUxTTmAmZ5K
G/WsT15xDR3sQdgfvqGMiFs/YCTZAwxxcpQmBhoxg4aRVN4hA0i6UmB3yCuAwTDtUiLps/FiSCIF
aAg9lqbqpvBcf4bQDLR/7DpxVGp5MH/96ueAq9ubtnaWyvXYsFky4Opg/sXwg/PlTJ5YLLbA3a/m
9dVIWBZenDDA3HLD2VqJDv7A/+yWyIkXFpwpaRM2ZiqBg7sWUoIcEeWQYeU9esK1rKR0venoMCYx
k6Ebj8SlVIEu9nxKfVp3L2JVEAyhawsKkrkc0rAfDBg/xdhb54RpvVKBejCAnFpiS2dnzSd3IgjL
DZcjNdrq5AboeQgbmfw5RcHf4DOEsxC+E2RDIo+r1+7Dy12uUcR8TIY+W3FDBX9NWteDGaWjhnkM
Qub/fLbM6C3CdoSGszD30C2h7+2ZNSKr5VpMjb/1/TbEiHUnYS5LCM/LKIGCYXyh6wgCNClfIjQH
bPLvxSmE3e9/uYQL1wLq0LbBeHHoDtwypxCE4VMtp/Akl1xEo8ARzI4LUTxCrrodSjxyb5ymrAr1
KRQA4vV7xMhG7/FPiCwxiK3wg2cub7tojT+MLSfgSUmFdUTIcKwmD88T6j8Dipm+li+Q4bGLrGcW
LCw3yURYXBNLwsMXR7rfJMzMZ69C/OriVo17MP8BAPbZskzRSXQPSYTr1A+1y+INDD3YgpFoGbmy
1Tj+hni4uHTun5TI/41Q4oXUR2jmnRMTWdShSXMJa+DPyrM0y7w6i/nFNGV4II7VuX3B4s1Qvokw
nhBOnW+BcOp1GopN7yJuJirIgRK5eXEBXkCuU+CH0wpT1cQ7BKAcTX3CKdZWQGP9o7H1b8yUsxYd
jApF9Ic4XkYHN9xmGw56vxAaDlLxOynfJ9H00YGHQNGC2ZEFrgrqBgNpXwDNArrA7Ai9GAr8B++a
RGhZi0gB7GeKjSWOeY8vOC6ir25dAXFp9kp5yUgzy5L6AYjwPAOMmCmm2wdC0ZBjzRw95vHj1S/Q
62xizl0VQIwS8Xvq7zeUHuQ0za/RUXjmQZmw41EVKsf9KpchBKPPxKgJVBQ9irggbFPILGjcU+dg
WawDNH+KQqy7bSR2xNvHwuunefvnEDRsV202X0znjmbNmcGCbSflhRo1DQUgyzvTcx9uV/5B4Xkk
WamF92NhBhkVKWDzGhimgI+SKhZF0Fn9OY2JQSesxhwYZkQWZx9bh8g5eryQKhVEh0IaHg4BG1E+
fnWnYGn20R36XWHGUbmoz2gZ7xvLEKrY4KIwCqmqEg24XQU5WFzvk3HSIhWqT9qM1vqJ8f5jv/xI
9WIKR64+nIAdIUb729z6pLo1+P24ToKJEO0p1n/yh7QpQ7GFtt3jcaHMXXg4jrm85ufKgI4iVuDG
HeFnS0KP7Xxd37o7KRIbFErQzK7OT/utSBdgU7fFBGYegBkMMnkGkExJCOkY+OUVe5piB7aqoAf6
JsYEpoA/9/XjEI3YVx+wjRB+rmx7ikQfd7zvD/Mu5HPYN/6/jdqurFuwvurmrwNxnjxPFBN/zoMP
Gez473x2L4EG4AzbNKLJ+5KsEQx5AfOj6cYoeziIjjTvOYVz5Izts6iNfC11CTzZgiYqf/DqQRPq
1SazvgB0rq0BsGu5zM6Z4Qre8UXjEVSwLQImThDFtjdUYhX5d3vQMfZp7QOSMi+hgF24BDPN5AcS
svP0/Ifj2N4fjRLxnWrTUE5ZzjIRJ4tG21cDABmYHKy/F9ACBxyR66gKpyMGMG9Ojr4TXJYvM3rs
7P0ZpIPsaqKI9Eki8a+2CXjFJeg7Isowsb4bNrPwY3vUvcrFvbnCV7e1WAF4lVBkbvzqPkadQVh0
TeDDXxXbhOA5fRu1UkfYfiadait4WTG2sP6tw0NYhlahdJ+BccRhtGs6lEJlvLT4gBTXp+Jmxjx4
MiFzBHWeYQ+5qs76v+wvPVQfK4Ayv2I29JtfQ8cwLJRm/LpUESy/Bbs1L6VJx3f+UaXQP3mU6Gwj
LM8/KutaYfXSbrAtXHGI8T5OVaFoSH/0ihuYKVbMJyuiveBo9NxmqrYn6eYK810IrQluwXUhmpgI
gtWUYJQpgERl76WXNEzpP1Rw5Xc2R99IijyB4k25PaIEcb9c9ldgrDYYb5RViG61E1htXp4N9hj7
dj+ZiWsltaTUmWXdDhXHy0I3ekOb3o0TQ85FxX/W7TjLS06Ewkx7H3vexTkQFtkQ1pg/8Y7lfCFL
nIiVjVS3ppPkvUEW6k+EeunTwON7ffuoTBF7ga+Z2iKVhPBSy+0bg2ET8W97+WIseRRv/UPiR6l3
tCTlH9IbS1Ez1jygcFALDGMicuU1Ry2TlsSxGgnq66GZrXZ/2MU8O2DEi7FuZdRgR4FICTIhtdQ4
c2Yalkrd0jZIjL42Wm0myXZI8LvvgH/khznugu0Xy6xB/pG5FOyJeSViaU7YxVavixsfkG11cMhQ
iQc3LN+mWnlFmOuAdpUxB0WE498lYJQNWnA6yoI/6HepmDcOovTi8FsIqh4vODKISE7hcQV4jRiw
O50qaYdaCjbDTkZNuwubJIhwBWvGFqvcz1YfQVDsAHhxobTeFrJBvuF70C9/TIRl4ZTkvv2IRU3B
FALZ4kehdwlXfcML/bMA1nTyAPpyVNyTax9jbDWNdEJt0oE+r6EOsCBHJDj6cnjqdHWzeNVFoNcH
HD7HVOmDjkT3owpxTZfHOT67pHD35PSjilnuMQvgJTqrRxt6lhIbYHW/A6aZVwfRH4CUJL+bdyC2
0GdLtXNFSXjmFItNH0jAA6BjI2+J7DgIGyN7Jv+/GS+iuekZbto1BLyJbIaeYUwy8YjzZBZ9WT1F
KX2Jc4ZylfI+tf/fRLu+BS+Ms3QzyrSiqNFnZm65UAaB1IO5TMZ4gEmcfVrygMYv6oi37JRjxsdG
WIEZOB7luKow6QW+sYa1A+Yrqby0vc9+q7pnL1PX8119nK/DMKwqbHed6OO/Kz7ShMPLriAh/tgr
grzUg8Nc9+3kcJ8x5u0BNfv1ZgtKoGTJksv8kMv5NJE+GI60NSVzfHkQBo3/5yYXiZ9q18+c4TZ+
yMfRah1Btcb4lNN4o6qsDQldwXHdo0CL7nUjt8RGCV7cDJVLnus327OIrR2nq0NlG5C5WtmU8kZ4
GRjJKOeM7qaIWRNd4S82+vPo5w4aUPTcD5znyLY87cyPT9Koh6qzTI5skMLQHiEzoAtiEsuinvw8
hI4yCXtsR7UNWBdAOFX+Zi6iJRSjEpIVXNkXObJ0/R4iskcayMFageiEplypSB3wL5Xnh7PG5bd2
BQnxnv2675uJetEokl2z/GcfZzbbcbwFgJZI9DiYfY7gREZ6NQR+kisI+VgFSEmmuuUVsUDhWWLl
kfa1Xi9NcxuLbVSqdjBsFkzWxdhKqZZj6OjX2fdsAAsLJg8CjaK1CoPRg2ZBVdLITiN9bKzM+aSG
J4xsUJVNRpXmmOCQ2IIRqGCLemTZ7Y1LNbHUNyYtN5kE3vkMs5/dB6MLjSMlynqjSdMXfvf+rZtM
MesJ8x+HtXx6DBAS/9OUH6z99j0ZsOCH6D04okbW38Ax7gyJqt8MwWtUQ/FNzrQhQEbhx8W90xrr
GI9GpYYFb0l1YDXUw4XKzCRnd1iebG2oK9NmsFFL4RRvevbBH5d15Lhu8jP9OD9dWZSRH5r5iLFz
wCVvQWj5qs1I9AndTfERm11mteRGREOFpe0ASr6k7eLdOzbzcbEnDlViDeu+wPse4/cKF35dc94I
5qttqLwfhF/GK+YL5OoiAAPhPO9B7dR1+58927lEnojFMz4tpHgh185IC6JjUWc9LAYxzNkhRntC
BbAyMAYn6E6T1RFrew0lbt8HTzKgLTkX1ID+u+iklOkZ0BziTdXMk/eMN+Nz2qeM4yljXCu6uSDF
f3f33vJhoyNjf25skfDgFrw11sh260JTGxLAsIpx3TJZYqo0mAC1clluT22G0hIVRTaXUQ/uR85X
S1ak5cKu+kJ/EaCQDGad7kP397poKH1Cgmjd2O0TYwjRDce4SwQJDOdl1CXwXYwEIGCmJAAgi96T
E5xisxh+F2wXBoDVq4n9uLR1GnP3KLC5tQoaXMSb8k7oLzwef7ZBwsJSEIuUaSZ/S4cacawdnwS5
VPei9jpmItPAUyHiuAEzjNBO+GsflhsD4mSxtESVgdDy1y9bTne77rggTwMMx+oukZ2DW3Yo/9Ab
ZrDhiokwjypMlLTr0/vvx5r1/JxTXFpDpAvZKuKFivRugHMrMHnGPDJCi/CIMHhj7vNA0/TQpZG8
h3iRmA+QsPoAR//SBczb3FGGhlZ8RNwVktJh9YoOKjnV2Soo/VBljm66iNp56Y0IeRgb2mENjPPV
Ocu7V/vpNzxDyrcMu2L/XEJrtGEhfS2Oo+/VsZytFoIxI55qFXZdyjrlMzLpHhT/BsE+VnC57LsI
wDExF0usC108yxa1iq4GEMeV6tL+qGf3cf+dtVo2Xnus2UhkwzuDai+KghPLiyG+r0ju8cOfWwvD
v37iT+LXOrJR19rf/1GMoIjWfpx/56LxRY5hWYXVmOyzsAdGeXYookqHwzMsg/gzpF1O0o4oF6LD
iYuMsA61o6W8Q+Hg1Ww3oFw4xSPPHLHGpFE8JeQ+7TF//t5o/Wel2HeNxnOK1hVvmI/yw19VTypU
1zIH9nXG+AnhqpBw5/3ELVbN3G30m+hs2KdFCh/TXcLo/9RZl5TwfdRTHlr6dsYFCUmVXl92RYZs
iK+V4fyafpxUBOX3hfvT28noPPnaHG8R9M7P6sqOQ5RdO1eep1yKJT4m/PQxc9GXTqMlZokXVO0X
K/TglDbCOk53Q6wSmmWHslNIIaLnCsrNCzFaeHPJOdp+/xerBEDJHlYoeUYmoIuEasfhUQ7m6NBG
gQMPe9Asa2s0kf4r5Etmq20ylPqzye6x7a0JrAlD46//rUfQ2lHcBK7bmAdGNQ1EzH+11lEoMb0J
DZbngmQavFPY6EUtXSonaeullnbquUF3VGXtfvCgTEbcaON9iiePjeViHJ3r+ohA0wVouwz1kLJQ
GTE26jAUdW6yELrisBMMwZo42fbeVCE96DvXm32jLQZOplTVyzBj/gTbDROY+7A8SDl/5ra9Ad+d
wkx01uupuHQ03mb8KkEQsfHxwo0MqzMvhbEWhTBCsjo6VZleBzQ2tJQxuvzthF21w7gVXKyEXKtM
3CciV+o8oh8K7S6ctBIueSDdS7jZ/ddwK7E5XbILwKbYquwekgblZzsKa+bhE1JtIfQMsf+xyFju
bePA03Tk+UCZf6SbsUEOVCWBOTHa6qqmPfY9KBFh95UsaVd66ENUM4JPaNvf6GyYAxc3pc7CSlC8
20/Lf/k/6pn8vFiYyvGWgTYKCITA3NolGxP5NGShC3m1lwPscQs7LIySA5xOVUk0GX+jzzO/3LBo
dnSSAwS2WKt6sah3dBqkyNpVDiMYYXoK9ZzdvyIM+2lwoLuO2jpDX4pXCKU8PNFzeCuLXLKRt+H0
PyXcUotDSIxAxq9DNam3Wm7zU1l3RKQNtA2ohOtCVdZeqW4lyd0Uwuq0UrH3T6/hYSwAsJf0l98a
CnBNCovvweRcOvrm/6/20DsstKbkbhPmqsYn4EXYpvMWrqYogG7hjU0bqIbYRvz3TqzQKeL2BJm0
UmjLXQXgu0YyROvoPSPHa55E/zlfS4vAuURq/YZ3EkI4xii6M20Rn3pYHS3HteHQHRs/5A3jGMP/
AaCCuG2Ye0Idk91VFA+bekc5dbfctTlX9cQb1+dy+wZGFDh0Tt1A04D7gewhWJ+4N3N2U21lZvYu
Sf0BRU3UttLh6M316UzLF3m/AvZT1wdhubYmzvrNMom4Xg/LrkOPL1PgfZG1G91oqwnSWykCeIQ2
+ctNR7PItXm5NFmPugYV4ffj1SveVrjseUMX5IslxPpfo7PYce0Nf1NAHsALo5h8bBlkhdvhq6gP
hcYfyNk7KKeSI3H60t+eWdUHr1LLU/EKYSY7HtiOBP6+IZ1SaNDriAs2mO0W7SKyLvXWFWQ+lb+4
nWDGBDdmBRe/QVZDCXdFSrxVD62XMyyweiqYQE85hH1P2xbHMLuP0S3mC+qMDhNxG5km7OWTbmI8
yy6nHDjZzXZ8ogO8+a2gwA+bqXyhuYlMnwEEYhSWvXA+p1mYWk/jwEOJKUuYjMjyAo4ew4OGMPBD
YtxQk/YORN/vzMbE2daqT1vWbkc6SDFQS/qiFnXgm9jeM5+dPRuPEtwyXAcZJUEwfVsFtpcPAiO0
VhTkEnfC0bK7ChKlRAb6mSOWow2cc+tkK+Q8prNkCJrj5NPLSM8bCUn+Pm7yPIrnUvieoBAVZQKw
R/MIyw+WhzJRUnlPQmtv5A+pfK6RbbV5YU+82lJUTW98SiskNYjhOysauW0STpFPBovq8yCIQ/Ok
7O+cwHvz7STyMKkDFQJo5zF6I2mYVcNul8MVPqrSxlt15//Xu9t+dTwiGbDzTQFPh1mDT/61O5AJ
Ar483FQQnjnG/aTz1a4sfcyh0eaKh9smIKPkuZUCjUKPRnDKDxOV8wxdzE5e29L7LPk9voKqBV4t
PZZXyNYVPcaLHYqL8zbJi1jkMLcOXV9p/HSxPp8DWxmK3ABp6n9lrci3ip2MHOfuFe3pgMRuPsk+
0IALbOkfUNVBLJIP8/lD4eSBTbdKoNRqUrpvTcNQs7Uucc0Y3CZibwILbdshbvJTl8VtOQI1dP62
puJmjxdfDja5iSMsRlxrwPWqkyKY1RQOyXJVtmlZ1JWxX32NB0g6hvvRl5C+hRVp8Uor8jcA6Ozl
AYPrJLotYStdI64CT8fNlZL9/IPKAczdDkIixhhyTTMuF2kJ/2rBYjxBnrzOfedtD6OGx0wf1VYy
wTpiYWkiuXDEeyxQgEEA2z2ZBtvwwdM7AI1D05Sin50/vTRbE98+UvpnE/g4TDpB6Csc5IM85l4F
jRNcWhQcY+RQduJjpqnXXQ5K6T7vL9+pLuInO61CP1r3eZ/sQ6cSPMU/2sQSnAkpNpTI6x3joSPY
zdA97LPlKOxTieeu8Zd++BhYWPyBpvbWzfHoHLM4gUs69tW5wuar/HsGJs1cvi9pGGqSrwM4Lnwt
n/8ABwWKdcEwk8VDLIWLWsElaKeih0owDSwdmV9ykvNYviOIwRmsv8m4KCdSlvV782JngR7xVSHL
j/3tGvEhz/gvSjnoYlVjD0Q7Sj6yAT4wlbq1ERpQQgBpMx5ee2yzY464h6MreU422KlRFiEvjLCS
eGyz6GEbu0boAVGmJ/mcBLa6i+kTAFbOI2EURB3e+bN2DMvT4QJeK1iTADONzwAmKd9uq/Pf0k1S
0KAlWiR/qg8/OPYXlpFJER1drmAYLA/P784ZAHkHPqY0g3/pvqWvW3fI1zFvrgbExkJwhyvp/TFa
LGvOysX/Mfp3MNRARdsh/W2Eo2dVxueM+SFBtDjY0nJUomFrR4GOVmYOt84o6oF3dRUGbRqLQsba
K3RVnSBd/nZKHR9MZ9ptSA7MI0vu4z4xmPeT4dvlFxKy2iZ2vbiZdoBzuYLbDZIlctCiJcsokSOG
sZXvdNArop0MsWGG2NHIzrHvCCOHhW4EC8TAibgl7rLnVgZtHk+RSy5/0iJAl8EMBEjVJls9H/Bs
QE8pKs23sCc+TlBbHFYuZE72gM0P60iEMM8O126qq1h8PBVf5qntMgRL9BxLxfeyGjoEMNgglPTl
a4v/1HzmLDVNsIO10k3WAwByRmresM0egYkiwKYbjGMSxv0TU33VrZsMTYyymcU+IwwwoROamgE+
bWVXIPMADxqE+7PWKyXsPD0y8/gUJQJI1IEbPCfHziOWR5GOAkXdVCiS45MLZW3EInptmJPzbtWz
N4XDIRI6B34a9O7DZlGTLoFBL3sNbO8slCOUMfL7o+T6N0WQT6RAL0Hi0VNVeQQeJffhmknl/4PT
x8zVDA80KLZbVgZqumulxJCDyXTO5VMvDe1kjsIB0h4lAlE76oS2CrQMx7leRSoO+yee1CF+zRob
4S7d5YbsmtTNTDF3CtQ2zgrWcUeikye048xN2e8cZWIr2UaDtU3LAgHEb0oX2DZeMSGd8qGjbvOz
5PG7NWS41vsYxYbp/lIEh/7/7cN4SQl/9BdDcC2PwX0F8DxkknKzg0wI/39h7tlo5MeoYuL/qIh4
G4MoGy6/YZk2i3Eiz5HBIu/dAE2GBGyNzjM6C5IRrf92EelN8NqVND1OoAWFNshSHKuAA5kpvbyW
J1fO8pz96M+FTxsCapjxxNHufHG8Xq3Dq7athsOyyE7MHVN8g9BAYwx+q5ry8x5Sd54QqsY4bx/O
KgMJzQ07oE5Bo2Ziqm9NFs+sgZm05i8krjgOHCEOB71s0DGZ9/E/aIo8C0SXJqaXedjgGiFHvM4y
iGTmcT3vi7Lg98CTNnz/Rf7mklC7peBlvs3mmySC94gBIva8lJ5iHb8JqEWrMCor/kzSsS1vigrp
uxd2Vew4OglanEtTsci1laokaIt9xOlXmWxlV5B4xJonk/SsEUGRPRafhcoFXjlEdNFS5fNe4H4u
5lbd6smWgl/z442RisRvZ4gjh04XbXTG7gEqjPKBQsyQ3PqFULXRiE+gh7Jq5O5pFwA3nkSmdA9r
HSJVJN1gdQ7iVbltsmRO7SHHX0coSK+2eBcKzGo/Olxa1MkhlNzJoZ7HHwAoKQURfTGAK5l85fae
oiIb4sUBLMK0JCz6YBOu5rk/6ocLGUcuW0WG1cNd+zRSyO2z3i9jsIYLkXPiDIVhEWDcEneEDDzI
YbzkiHXlQxTpXIcgLqo94ZtZJkf38Gd0flZl0bPCnhPUeIOsb7kSuy1FaUO00RCqWLmFQvhesFqv
kJpNV2cvMg88d9agph57cSO2c9fMFzW3zuNljHjMm3BY8iH2dyObSEAhZsf+0B93m9h17KifCowy
t1PkTwGJLuBxjoY4krBF6EXkH6XoBohrLSg+dPEME0eWrUoFLAjQHQYtAI22XbnP8DiyYvhcoKVX
rrrzciaoWV1fPzCPkvsYe3nDA9LG5bIwgBAM6mP19T2KjJQU6bwX2ytGxiM/7Rr7XOjB043+suAF
cKHlCSfbsagUhCi6O5OKZSsT1O6LN1dPprasj2x67C2S4hR/cSQlMz4rx9x9TB9o7Z90afyHpuSM
dwFtHGUucfOFbgLQlnwD5GXl8u7CVsiDYLEuOZZs0GaRWaViuGetMAx2/fBS0jVXH1gZise0aXDP
cnGcbhai0XpgG3KY+rT/6WGOYOXRDY+hmbKG2HgGwoDK8n5BX8F6Z25UOUhIShbFjhFauaLxOh4G
eCKX6nRRnviFBSIN4EMy6goc/GHWE5Ah4g5Azrx4jqfGSeWPHYLuXsc8CLC5/gtzTBwFIvx53CKm
5v3jH9nTgcH4zCqgRO6xGktmWUyLucAb4Y3JBJFhm/LCdRkt/1/i8g9nXfRtwRDmrpCwfIvRZ6s2
RHwW2xPBaPO+U6GOJ0tnCTfCDXjijK1PVpyG5tt7JxKfqm8QG57u5k5Ywz/Yt9YySAQt67apEUeJ
LMCHiF5J+M4LMo+nSzZe/C8sI30bHYRbxXPB48nSK4NAdmqHrq8bwJtHqAtNhGj9HBl2GjWZgw03
jo4Jnl4V381IHHwOCDklEjHN1zAqEhxvPtOR3T0dbycilu7KOPy5Zla467nFhBjWlnTT8BpqY9YF
zkfGV/TJSpjFUgrDUC6+4rEekQSRdkJllZCQHFumAt/hDNioz70J/2VfCWLyZFvCQUqn96ZxmTh6
DOhI/rqvJp44RQA+jXtKy03KYtD6AAjMHZzztc1Pod4yCtBYAeo/OPeTEphGTd5p5PLWMwOQ3O9D
PClzlk8HtWQXJ3sjzI9wVnGHLjkdjzW1n+DghguFqAt1RSpph+kya90tWpoeZsXxbg3Q7g94ZFFA
bCleXpa2jPYXQHy4IoJ6OClpaIDjhJWiIPwMKm/4PtgO0WTU/UY5R440b205dXQLB5T1lliFasUb
Ql5ar+vq90kHmxDESIbAPpNCBrK3Qf59oAhD2B4YsTn8hFPfVHHW8vgvdneuuI5AsoxyEePiuGi2
F99H0UuDRkf7Ba6BLW6xWgCpMgBIVmaJdqnqq6WyMzLTJFF3HQI5462a5lSBnkqYPcASbuDgfMhK
SnyIyPv0jOMUPdPRf30j3OLOGLJN682vldGMWFTeuf8JogjUdX62TtzML51btmvNHz8ar7CPzBuz
cCuIlyI8x6iJhouh6gBhE6QuR9kzyY5EnYvxBWrb2wvv7rNdlVdJx1i6Qrim1R+t+M4cFhwzZP3Z
3XPEFzo6BSZbXVfgJvOh+xPdB7+fYzKbyhAFXLV8vvuRRkNFny/9GbjLvYtz3DcuAFa4u0EzTyBs
s1DwzOGIyNdUHfQMpzRVQhNci/6XaRdWa81kG83d7QgTB4JBSSab80ku5DSPMlvd4rbYcCqNsMYw
6NOHFW3zJXwsSPGKw1LVOTKPW3IBsYC7DA9UkHTTc28T6MpknnfTPQrM317/AGfhl3BR/92VMCUy
e7YK3VJ3WK8Hq/rAKEJbAXY3mT+UUKOWg1ryOT9xS4LAfGjCF1JqtYtHg7Xr+iTDWNmFB7Vq9as+
h08rZkb2eb59ts/FEkNMGN4gO9AYfd1PAetYCpqQzGERxgzs7c86G6QTRoh1y4xsBwYr4T5MARwM
FbIwpBhPzOfAsMjbh8LXemD+kGVj7bJzDsOdAqCa7aLZMp3ZPqi9E+EdWLpL/74swonj2LSSzQNj
DtyOtt5B/i35qKdaYTK7YuQ1rlUtSmY85S31nl5pQvDN+GPADeIE4OSwZPt1FPcUW/ZC+zYuN6XF
lpk3937Gw1dA0wxQRjZsIDLZR2FX9zG5DAFt/9bU7LAY2zbWOnr9NTDZa14LvAx9WxMcUF6Pnv0m
yySSOLsCY/0vsGRkXSr7sjfPeSV/cFaRABM8WHn4O6Da40gL9+0eCf/l+InAhtt7PRhi2kaFLo9u
VtXkpyJ0Xh+OA7fLIUFJ3IPl2pGXVfj2NIyfRDPrSHFdOM77T1edae1TdvQFwCNeaE17TtnFLvIN
zZKNMqTDuFUJI28VTPK0gjtezr8xiUyWPLD62j/18qMGHjwXXqS5W/mR7doSbOJ8gaPosIPTWsyZ
WUc+ZTqOkV3FcNKpXfaTx3Ey194PWQcS2+wkMfbnOp9Fu72LvxiqhxrlIL+sFMUiwTovokOM40an
474He3ohIhspALbK6dzaYWIm6QdXrjkYrqOeyooNWJ+dMA6/6OCisx5lhsRDWT/SL/9iBcrgUm3n
T/LB/PZfXguAhr7JbqBbDA34iGAHekCPrVWQPh/oACSrEvmnL3rSioOWEEVx8+R6gm32Klcl8DZo
OPojfArRSyY0DpGEZqzRwDtrj2eauqBZFuHH5b9vae2U3T30CXh5E7YgQFY4XLLg6hSNBb9S2Onh
HoLB6fKkWgXAmG9ktBOZvRUVDutDVmvDWz5dNNib90Zq1flTAsUmDBklf87tV85a1ds99LbgEZV4
qacRnsTIRd3Bw5Ah8bRj8QwedZZY5wNz+s+rlMg5cbcVYqY5U2irz9sX5+nvcDHXzobQ27mM6ro9
AkeLGh/m2GEIEmL/R2v2+Ije0sy/BrysyHgDVE5MDpwtWqAy+WgBVAu0sb6xxup8nckIq9ACagC2
C5X4UliAz59/Mpe0KXU7pc414U4ZwM6Uh9rHDWA+Hha7W8E9KYNyRcEgIuyiPAvzxkJJL0kVNYr9
eLDUG5h4hHQg/ogi4ZHoFA46p8B0bwaMxjFuzVQVfNECpn22VyLgRpz1rALQlvRAhBdXVKC21Rqx
X2WeinaBoLKIMD0Pjc26mcalS0N+HiiIX3WbkGIMgilhWRvVFaxC1/soWlb1J27kkY5WMjeQ1LsW
HM9EwPsWeGnu8GteaPuq/FGwZXo0PGz1VO/k9IMB/Qr67qJ1NXQodmoqvcpig/Iv7KrJxf7KdBJU
fMCc29HZuKdJKTCv5xv9uuZYQqrcWowTHBcwKmmcEH6BeH6DPxTjW3ozU6rNUoQLpjla93VEQ/T1
Mlke1m1FtUofeJr+2vTLvduzb32qklMrDFlgcLP66HUeQhViAe90G7tzv3FpgjWBQ7Gjg97T294U
EF1zyqouQzE8wX7n0b5+XLNC2DEGEjS5vCDdeOCbW4MjAIPKkOTKVxC+M8Vvi1UrgaNkkdixFcoK
TDIsHwmcYM26y1es/BBzpBXZJyplYFTRDA1P0b0x8HEz/1BkSrHjOtTNFfv8pypVrIx1nTf7NT3A
TuvFG9p8SPxkkj8YozDayvENqzdUCbdtS94it60YttiXtQZNZHfaPNryRKCgbeByVySqnk7CA/Cf
T5o1qXm98zBIoWE0b80wjlZkLFKABw0GW89bEjavfI9mqB9z9UtyBlne37SxyRcnafFfbgm5vF54
1l/NvRvih7x5S267oAzW3nyWCJ9qJWqh822gAMAbwHquI/qS+bIL+cJ7Al4zapjhmDI3WdCrxkEe
Ev0TI+B6UsB5TozrECrVtvAMP0eSD/Cg3rfC5l3PE8goKTlxhO4bvRRMspPx5TarcPsijbcqqAvh
wxk1zyHd21F+jQ4L1DRhq0pinG16nJZB7/huQLqsNwT5f04fjDOwRDNBYL5fKXHI4DJXrgu7m+3N
IIbZec3LuFuGW4ld57fuqoW2Jprcm6Aot1quXnyilBqZcZeeZTSKZ0QEg0ZagXCSDwTvqTMchJQv
Jgv9A0JeuwQUHk1Rldo/NmoNO4qML4BUT22gEwS0+oVogsAjKAxAeRSN51set/Om3610MFT384DF
vyTTBdastkNrE+yfvEt+xilMIBMpRFKhk8hWd9n3KEblK9ib0A+7jb17tGI5og2ThbKfQ+EkGuV7
dQXhX9LdKF+rp/n3pRLfzkgn+gP5cMllXzRtGwSjbS+CFOWfKDwBxd0fA4o73mQUNnxoXyfu1zWG
cdesJvCrwPDKyH7jAvsxhz0oEx5+DAQKjNul2KYosSvjqndNiE4KzFajZLVqhYFivTw04DaQFP0W
ooOBjjG/EOgZsU8jTtWpY77Hq/Lf6yFCqRl277FdLAKLxQaJghQEZf5OIAeUi0e6cQ0iSso7EiCC
YI7vXFvrq99YYHd57aIVHgDoI5r0UmRZ36kljBD7mzkaZ/EjUHTpG9LzdtqzX00P0XgKc/gM8kJT
IFLZo0BvzgXTih2QjrLMXvCAVjG+Hh5Ml26k0oyCU9nm3E6XNRwwiHblgGhKaOJAkYo6odLcRiKo
yrnCjz6rEjzXFKeDZGrKKA/mJ7ld28885W2mt1zqppC1ZxGYfCerSDMxs2vO1t3TL6clR64MWSaK
KM+iiikRowFdKyxter1IdlBZ4oJAEz0fHWyhu9eIuxKVc29dUCJdNiXH+rEWojyg4XzQZ/Fh2IMc
hs662AXyn7t+SjqcVShHkqIO9qfE5Mb6PaqhAsoCUz0UwdqcYkfqe+xPTkIl8vRdaFCB42VVIyZV
XQjRgg0u0N1OSmenquhCOVatWCM4mU9wa702GSTYF+udgrqDMeYwvgz+prgFu43Uq2ksth6PIhcS
DSnNi37aoXdH0ie7RzshQodztm1EwDvHu808xNcbGaAA5D/MSJQI67LKShG5DVaPViKGwLO6PcEf
abF611z7JGcYn+4vNyoEjmpdXhSJmneeMhpUe86zpl7cqfTFUYz12djEvrzJCsyI6DkzT47DtJw0
LRhPr0ZNXxXx7hsyeiTQO6u6YyOd2bJrXW1eKzvWJIuswzqS4tT0n9fBYMvmmkMOl08df5cfIcsY
rUpl24KF/seeuJ5kDeOHLHKrYDwBAhQ5tIPKNPo9c/ealm/uWTf+l6CncYsoOK4I8irUrXY0kOp+
3CDny4ARr2bFHRc1WA3eJqS0o7BvBCFMtfYKoNKz2mHvXiysgSwUPx35ZE4NQDCxYJ+7ywAHOwhM
K8WeyWeXDedJJ7mWXMC4ZqPnoKhN1ut1Kxqj2E9k8tf4kyr5kkpRt6CTYYI+d9mBcCsn/SUl9mEd
1wH4lz26VpUYgPZSduS+GS8JQ3zCJ6ppxhsnB+4UiaD+7COCA1tpwuvPunfLsIyUSbd8iRWwpc25
kQ83BtZQ3m4LjcEGfcyeV8X0qyCxQSATQB1HiLD8ktQU5pLt5V/NGZWh+SWPUvTB7Srb2Y2lRFQC
tSGVh0WhSelS+3lmZrkKb3ixS4y91EvTbHGqGqvbFLEFIQl0SANXGqHtgf8ZrKG2JZ9j1EPtXx3I
v9SmeNshPwrtlr3jHyha+KU8CTK97QEFtH9trI/IscCKx2VpmDpI4VgXHuN5oKJ2lYYyl2GrTEWL
+xPeQGlUWXc/MNj/qd4huLAAKoeRL4AvUDPww+1HwCLFKnqvaM/kcsRxXn5+E74D2d5foaLJQW8Y
hzD7taXo9RNypNreu+1WjOjfuMP1PBpmwOU03rUMPpfPSLK+IAEpD9vSFX6NGx7ci0IxfP6mQJZE
+JQNB1a7wULLHexaq8b8Dwtoba0vsFEc44ljhe8+IpaTFMHPhxiIVklFMa1qqDzOwGBwb7pcKsBf
ZN4GpsGO1f5HwgYAeHWOVl/z/GKa1q5DvyHuPYHBse+eyIPWwt9+z4EoXXLk8VadcWlZmIMwnDpL
kFcGPo1n1Ell2T09tXcAlwFWkTdD6lrnpRy75yTTehj7Sd55Az9cbwyGvz/InhwEhJRYzLPbfduv
XOPGfUAWhb1yZIbh25o/MZvHV1lKhWdONOjjHfdI3zDaU/1aRLmiQsz85ydFFv8u/PqRDiJX/nwg
ZDbR2pQsXjHFYvdxT87q1toa3QIxKL8U2cngqgaFBSdc/6rWMSbrbVZu+a7LpkzPqR4aeyieMlO9
v/G77uy/rHQstC7V2GiLbSGzJ8cjiXuMbfNa9lRgBtQ45XI+cwfdt/X5qsLCRN1IZg9o5Lm5XEeF
OP5qriCupWlOHZbGRTxHCwCzQ55KrNRcpIqcLSo/UqcRjh6enWmTZ/k2Z6LPkTezMlF2jy1i49ME
MiapkmWd2y7UeZy5Oc2r3bRwtJb0wfdFDAffuf3GlYW0dRnx/MDEXz0HL/gyiuqy6E04AXSeNxRe
nKsLxtQJWxOb+rdtTTfwXqtafFmjCDury6mmgpms+ls2AfP1TT/DJbPLcTnPxpVsGUd282sq3ltQ
BbmViLuKCn82FSfMyQ/SzAbfp2JkVupwgJogajkRXHk4TRuUmwVNqmB0Ogw3PwTPOND8QusIiHwV
LwS0WtC2KBd/3gLWwh8hVw1fSzK77Ymahe74ytcQyN9vPiNGyG/IX9cIXkFAtewAQho05uQ+YcBv
1PmlifFxnASnUguZ8+lLbK47nFnBohUyWzHkMlznyR70Bu5ncbVQUnPeYqLP6QLpPQVXMS+Dm/V7
64JlweANjeirpdqHHxXx0aWh2ql/NY3zOU0QoUkdvyVKwJDBn0EoduEUGlRdTxncoHahFXAwfFnh
FhEXpLPyCeLkKdZOBk0mRh0AXVQQqpOB6Noew2AX8iUaWqIqwawZrmVsY5tOWbtAu7MWCgIThO/k
AP038msReHFJxY/0xx8F/MyXq0tqGrAyEBV3LVaz7hSyLUsTRR46X0ORXL2X8VQqGK8CC6aErXm2
BcrY0WLaOL0alfsRv/46j6OZsYBODOIhVki2fVFPqW82NrsubMwHhZ0xtXExS1PT7prmfV2yZ9T8
AAPQyl4hO8LV8+h8JljnA4z42/Q4jW5z+NstEVLokHe7L31NQNEx3WGXBcn5QFqSpLseyEdexGKb
YCTA57zRI015PSG14xiwbNDDzqJzDVHNWoDRWRtOqPM827YoGC+DzxGGgwKMPs3obVOeywd62812
AWbLfXpakC+zzXdtrWRCp9Zf478yl118oCOQ8Djj+wBQGtzlOFHTUEUlVd5qv8Jvtwsq1zG28/qP
M7fx8C99rOw6mBusZkpeuyxc4QkpW7Z6F2oI5kbnKg6yMUXwVlqLND6RBQnS3bHCf6oNsPBCbo9m
2DemtJ4Wha9eXYY871v1JvlBJdIp7QxsHpmQrLRDoIXFHLPqB/SmUAxhYhTaz1X1LINeSBTKqHS2
+4f8Zl5yFa7OybF6Q+cp3KsfTECYc/0U2UdOyyBeaau3BrnV9/xfaN6kNfJslnv+1FmOVH0M/+e9
qdNQJw+BrWDyVEtvzcnFHNHYPiFFaA/pyZZRnnqco2sMLoJzUYroX1mlFekRyFoEgDAA9hlvb1wA
DMiDCz2ig9A+0NnaKExdDsH+njrG+bXGhYPXFd/VJbjkUMeCBBdNSDBFPdjGiXyc9JlGM6BKPQ7s
llgGAeLFN6NzyM221fylNgk93KRTowuEW1eRQ3Hg+tM7+5jHJVgGlX2HUliEO9bUVVZmWY+Ql/dP
uN+evHIrMW1/HpjNnwNzgW5aMGS31A9WkTwB803QeNzExQ0NdGb2c1QN0LfoPX0op4YZ3OEbXCnW
H8bvt1bSSFiM71wHEprkD9b1hAKA9qd1/x6ieMtdTeZImaSj3sJlLPvLSMG1QraBqPg/Bf7FfMpp
Zp9V2Yx3qn9QPoGN/n1mFMOKg9mh2HWXH/d/zSW7ek2zfjM/Fdme2sZAY1L0pwci17O1H0xXYaPb
OyN66Iv7b3brWYZrtAyX8IYl6ixxVu2YJf5o/GLUt6QiB2ro0aQ2lp9ihgpvKtr0Yk3BfenBGhmU
pBKg4Or6OIYzxbpQtHqSup8xP3ZYcJ7bf2v70Q0XKcdKa6RIhEwscei0/z0voyWI8ghfQ8y6LDHj
2VI80ZecSKtTK/noORPasfVmCGT+j8waZfzIVEt5SqolkfJSdTkLGy/u+VukpF7DH5IGY6bfhhTq
ThSfJJhWp4pcjw4PA7phyOcq9gdPvdoFIc5czfNCkmkrQiqxnBpt5wd7ZqVkedRiSoHV8DsR7TUn
ueV46IkvMuPbToyEWjFc/aO4MYTEAJezejv9gy3nvWPHkOUuVEX2qgCoq2qw4S/eIp/hsrC5q4Kr
A91FPVMwgj2xp8QHbsCP9jM9sCTaB4EcTkwTE6j4dae3BXEGJryJB0bGrdyKvVD3Gk45GlYiWsAb
8HWp0/TayXQWM1Px0Z1p3KRTb4w2H9i5zasbEr4zeQhUieIYCD6+8eIt6sFPZPvaZ4j8t0lvGawK
Yo4rA2n9hwXGhX01h+1ksWIH2jALE2j2c78XyNoEqW5NgO/CeIeTxn9d8cxuUdux6ISjXcgDTPAk
tTYfmsPEBgqnpqaLe0rYL+tVGXABfWMZ/TtgfAg+uVjgfx+lwyhNdfjB7Gkzhz0NvxnyaNK2tEl2
eHqF1IZMzVnaUqCAiptnAniqR+owpEFFAz3Mihfr1vOgCiNM53S5Z0w9KIP0cB1Cdn/jHV23XFeX
xSMcOcnRtRLxzy4ZnAFGZWaBIyCt4LQxv8MOStKXAJRKsUgCLdq3bK47IaXoXSFjHN/gi0v0G7aP
FJxehpXvdwnzGyj9Mc/QLD6i2rgPDjc7Y0ALmJE8oKbh5ntBqeE7draU4lfObJLcOYQbsxhsKMW+
xD3P/d53tKSipgDh5OknHRG9nsQJz6utfv/0xAi1v+NdFqWfrKKAdECWN2ZoU1cz91vOphl4OWqY
w3ncutXS0e0gxc3+zbFawY+bbl+xgkvBtdF4MRLVGGx1aZ2bN7sLqdl7RYKuaxBMC9QbCfThp/+W
R87lSbYK8YzQVfzGlPoLPj0ZzoiKi7AeE4hJtTeB9y7ITy+XPmbicOPrFO2X+pRsLSWEr3mEROFW
mC7DqzzHSCyQKGsGDXMfh44hU8O654y1rCab1CT+a8GhZpIfHLyzy8of0f4OOQTrhF8oYuX4v+Se
+z9zbUQOqdoK2RjxwKJdUgY4MjRUHF2XumKcp6WLFwgAKQKkAvw4VL0M2ZJ21p0noEqOLPtJkRs9
VE0c/lC2A9gLt0JhlLCaIbFR6SNaL0QFkcNTHnmn7eus/6W4K1qUEUdfk+Ejs9k9Hx4WjEGMVi85
bxb2wnHhm9RymUnjYFwPMa2+Qb4QpZEfezN/QM+yqPWNK9OMht4tsTfDZmWQN1FI+QZ4CmpxWuJW
30Lej4nOKNBs7nEi2vwwViG2Cl2uuijB2+eAvmEYB9V7Nuki6ld+dEwI9/WdFpm0eNc6M2FJlG3E
eEOUUnEtfciREMaYp7QpFhYoN9akM5S7U0lCurv2z+KoXuzEhRD23YMvkSCWFBn13b/EUZ7BYVi1
I5TztZX82dEp7r0zRMDYR9naajIm8DUu136kzM3QbQUZozCaSi5KGzJ0e5r0x00h5VEI6AOUdK6H
T2UHjZFZVDcjuAn3eKCWP5CUpifRoFDV7mIAXW2ITxvqwyQTct9Ykk/jpR2ORwXwK7lcga3h3TO9
gcc5hV6+jqLCuLyXxK+4qJcnFgnQ6kJ3AMRQM6rHGZquYKUWabr/yHaL15kWfpBUWq37KgC7rOs3
NxeeOPm6e0h/onZTf9RFwAZgqMOLtsTrN9vJZ3+sMpYM48oJjhT8PrMtWEyMfPtSi63S62BVdJtv
8+0LApyhuFjKPCC/NjoBlPvMarysN/kw4xHCATHJ+ALRYOdGGjm0NLokKwdr+UxC11cJ4twiY3Mo
Ll/1MbDHHacMgJ1fCRE0LQLYhQHsTzeaLFip/2fvC3ecyZZdvSoiEHNBWC/glyP3s19hHpbI6P5H
Me8rKy4Dn9z9Y/P1DUVZ+pleIMbDec62VoBwyA9vjKuOU5/5JtFtpywTRL0dA28kg6pvKnXcqTRU
0W4ndrrMCYJrzWO/9N0AStzzgtSHrwdbwy2yI4yAAi4rcNcc0GPHokIK0fZe/bT2VqBSXYPIQUGt
8H+6Y9c7Un90cW3+3DfbJI2i0MH5SWgeUVg5U1HWJ15QHpqcjLwB0f+lJVNEbeOeKyFmVDZwbpPG
Gs8rlx8X+4TttNcs2Q+lq6p5F+z95zdK2mgKhppXOhIQvCilhGhov5Gqt2RgiCpUs83j5DaZ8SQo
4fwifecGN1R+s4Zc2vMg/2UDqDTPbqAjD41gMu5AinJhyuM7u/McJuJ3p8ReUrq3y15eAqX5yBi+
zTAW6vlUi5KwbFcJB+5R2llJfS9J/zuNnjK9+LX2pjimIQqh6FeH35kKR6RklMQeaim0P6ivxejc
jXk1lYZod/rxz0XeEw3MgVDziF/0HLBsQV2hesq3pVHGMJoRCJUT3EyTteifPw6byD9AhVuqIVAT
bN2EGy06kO/2X6uHo0nMn1XZJ49F07rOD5FAs2eK32QTxTnr7cMbGqpYmPBIBQUZ8MaIKfdGURiY
TH/gSKnnt2xbL15vHgTLT1/+TCjm2rpNWRrWb+CZnhkqm6MyYlxBWtwnjYsFrGy252lE3hN6ExA0
4Yv2SEmjpV4+oatHUg37Z2jb/hzmnH74CPIyK32VVIF0EhpE4DpIPIjRSPgsvkEpCdyFddQ8Rdtb
ikbKWUR4hZdGplHaDGWIBbJS7MyQXKd60kDCO/HkL5LdASzxCFam90E2DW3l49rUywnfCbHZjWYV
H3O6vsUyVb8AjmWuVt602nyWt2VSYHjt12kmc3/ryzm48kYZBdOvgNdQP6LejAh0GHR0Hw+ocjLw
jh3+9fvI/Jb1lqXYiRA4iKgnVbB9e2up7ofgW8PYFatHP6P+lkgKQWlMQwZDI7cqJvW4ec1togoF
eK6s3Ri0RNDLsaoECdnU4k3B+6Az6pMmxfKc5Hy1DTlxQkmIfltgpvpMxps0srDgBG35dtDAUduk
dZTrfvQptZayyEflArp+nPTYomB27lY7LInSRyxGRTsYsonZL9ZCtZ8IUjzHjCw3ROS3wYOe+Myd
cwIm2yzYmxb3vTGsQzjhaRnnEjCHS/Yg9PQz6n2VS79Oq6DbFihfLCX3rfhbBwqHz2LWe6+tyLEg
kg8kif9DDwW0SJyTVZd3Ap+Y6PKn7uT0jJ+WxHdXP77UbbS95ANf0XNF0vKf7YxT+Wj+3A7uO1o6
48edoH82rvRGDjjTO0GwNHlhQIGdDfXMi2G13uTyYKhL9bA1pO3uzZ9wRv6BFg7a2r7a+Zs5I03k
pOTYPS2XXfdMUMKCjXu9zK5n9ZKrFmRgYcObMFgRkE3rdZC9WtEYo/i5czPNpZ4p/dwk5LNCkqtp
Xu1Eni9YbDPoyN2MS7hzu5bAQLrs4lQCGskOB7x/LqcAtbMwXgtaThuRV8ngQFRpDMyB6eDXD8aP
b0O0ckyTuqq3iJAM029tL6fD+CM/EI23jqKvHbkV3U5+S0DofI1Kz33KRr+RHt7HnF9SeOrlzkjM
Fgpm4OBVI0C1LjxreM+fbZY2N46E6EVO5889nVuX3EBtGMsXR1Q1mkuAHHDO3Ci7qT+Mn6w4KBUh
Rf2HUmVbOOIGVl04ytB3BOxIlqG96zPou4IKPbh7ThHvO5JVcAnTolEt/t2/YwG2BHJ2GcozQWn2
78ubaiiBeQUGFI6GK8ebdhTIsXHGAdoaIoOMuE2de6ioY4mCEuVCAcIijNgwO8DEg1jzUQS9ZpkR
VmZdwyYJcS8RF2Oboe4uvNyJw2LCJVqASu//fq8SoTPxmdRJXRdd/xmeMzcT/vYLALozGk1ocG4T
o442/oXp7rGJWhD0qs+0Ai3bFa3m5olz5CMEejECf0H8uZIZzGmdocBI54k/oGQ8HBZbRxD68jAL
2DGxNrVU9Jg4w15X76Gx+apl8pVzDkS59Mv7fagN1+bz8SCwsz4VCW7NB38PGaFjLVTQEqfFps3t
AOF7x82AbRzM7VLSeAosNch0U4K5mnbV5fZkgsJTDG6S0wK/o45EfBtsSa94wOvTsHo9rO6X4myL
a66i2JPLXweSFE0avEiBTwPPtybXzhzeBzZaON4EPGLNK4AT1pnXzAkwhn9YR3/PJUG7btjj2OEF
JcFFZgCUOuRm/of1sbC5xEcBCOwdHlP25cD6govUcz+SuEKFi5mX5Ak7A7YEhZHRt/bCG3nLBxgA
Nxc8isyF/aJG484b0jfbg6e6bqs3IaYUpBCTzJOffXp5326V0epbURUY6kZiky9T7/wn+QLJWg3H
Zwid7FnkkUxPDEGtt1uXuX0FAqCBAJpZijlDJE6Y1zwc6Xnt+NIzokg9x+adOHxM0/zfOs4TITyq
M4YW7JbEUlHd1YzBa9pf9qL3VxKidnsvBYGDKv7YfJQLbVrf6CPU0KCM5PrjwG1M4ULaBfylCK26
roBKvpPb/qv6fnci5NDY4aUr3H5sRE1EYsL4zITG7uJPGgt42q0D1Nw5LCcUJm/Qs42cDaW3K6yG
TDqqpafK/SqVA9KZqx9E497DurrymYhQFTKD0b7CnEMDSg34mZZrmwqwuYkLxPHliZHjIhvEN9Ve
6tPA6riLDRQXxLQMpltJMnnaBl+aHhaOx9HtLu4RCgE9ge2NDK7wmSePKFsJ31Nrn9YwPa5iAFO1
m+7ggsUjW37Pj31WszWTj1Cdhw36ZfaLeXUvj47VerPnBHbBqM7zcTEZiVj/NKk0F8IF+xWj5Srp
uB4jvMwuyVhIAwy8RXj6MKOgENoHovNObxbQ5k6hRQzxUnVGnuRLadYSYSqJvi80EvDJ1/qx9BKa
/1vPypy8qRuinEtmt+492RIMU78Lz90jN1+jCCkFVNHfIYKf17+x8DcB06o3zYVoQ6rw33uIbTM7
ugA6MQs79lW9tezfegOwgVJ0gKLKY3gsaw4Mr95hJ0NZ99eX5MyVpX7HnWsKtBNjCfcGbWBjAeOx
mBrBZlZvXnsMlwndDQ+/DucYoHI8f/n+f0jbd2t5x1f52enrvayrH1tNvK5wUiGSfSTvBg/1L3Wz
ryOFpxDOElQGg2muKob8TwnVbQUyKclCW4GgvroSch/07eXxg9RQB/j/aWt+ruuvrWdRk7Meck0R
M2n43iQ/wZk7+xW0zc9ZIP5ItvzVoFmOTLrXoOuAV6nG4GQgJDpEXcQHYeAmkthhFb/mQhQtcscd
nWwYeut8wf15hZLF4S0bkEmeCo+fZ3TO/rRUQBFB3XQ5YSHAVf/zX8Ru4OwDrWoqQ1M0JYXN226D
iuxRw8eZzB+QkUU+2PufZ0TIIUejUfpWaIdlC4j0DTR7NMs1xj2JAK/dTN8sXBJ7rsNg0w+Uy/8s
30oGAUkAHuJjP81uPtxnBqFxA8gBCuQMdGRvKuIhOIfc8p/y6FIl/GXnw8dynnMhKmArDSXYB+OC
I44v5djH3mUOPKSQYws912qwomiIMbwb6LmagKqCSwvUTculiUTxQQMBB30yOnS0qT4PAmty1+xu
QfYn7bFkMvULRhuQ4aUIA+2GIqJx8Bk7cdgvTiNDPq+ehlYFcGE8GiQtT8MgSALs8nDt7KoPIRrN
AjSwYULjLzUMOl6bxFCybRLP9Df4Cv1Bwkk8+CBo+Ws0ecrL/aXZIf+k7Byjf/YI7mRxD4WW9FGn
9oZVf43UXxvBGf1g326WR/kKAGP+dkyDTDEjIUkNLfkiluyB7eYTA4JDPsdrUBynmQt0TMlreZS+
aLla9nA7a7+PuoHIZ3sRY+dADOMx4/G1aiVuEP11qLtWiNWrCIBPMSO4nX4Xk/0IQpmhZTgXeIqF
bkMeeuJlRFvZPGzLEw8yuQ979/NLjgr/fXBwCYEwD0otU8pJQZ0q/SHFjZcAiz3PHzAPPDOIq6LV
4opMyJQzQ2vcvqhrJO4lVtw4+QWLtxYybC0ZzysT0rGT63g0vcAhsTl7+xiXjm13K6KPaCFI2Jo0
m9wqQ3j+IzEjeEvDz2f8H9SFMglpkIjn7CO3u1I5cU4PmajIvEYOtzRSs4OBjLpGB5smc7Th0TFF
ZDIMlfxJkWW4SH4RvkMfHRD9A+rrCALr/ardrrdp6L7wK0oD+PLww+ThNSjcCqMLaxYtsJdM1Gpv
tAlyMH75dzc7g1AdwDBsPTgdk1VHsjo4czAxU5ffMByvHYG1W6WP2lasEHsstkbczFshW+UEak5a
+4+U6xLe2HCC8no7eMe74Med4+AeL2arNYFKX1D9Da9zyhmBh2M7r6NXDu8bYwPN9tIglfFifxNC
T6N7xnHi6JYgkAtnnqeqN4yX/ubgt8Nwi0ubvbQo9HZFcoGE810fGFaoaXhNsuwj0MdkyyhfGnIw
/5K/avlmA+KP1sZ1EOtbs8FZx0QwNeXvPynBb0F7NxaiuAzLI2TGCIcIer+qW7fSpw5gXJH4ThZk
2ZKDfuAVOlYtC2SIRik9DKSFSUWOKLycblntxZFrrVTN6Fhw0WkmAjtLpcrGkXY8hogv0aQ5We09
/81eRVwnpz+EO3Wlsf98K0q22wcjR3LcZRBXVTYFOhp5NqjEpSIjTgUgWuaNdzLwqc0WkM0EkmZC
bXJ/TmCxP8xuh6fCjB9i9cF4Zsu5lgJ6CJKdkZWBF7fSUbWCyGE8aSDKYTQC3GytT/dCo/T5joLm
yoiMdgfj6/0HhT82Cr5iMxQ5hCWUuNgNSYNEVWJ9a3qu0xg0LdbaRllUhqwXB0qn/2qTrzIc1rZM
HXCcQP6HcnjDMpcgS70RrfX5QBDNLWglqCxfZsoh0z/+nbDM8ajX53c4G8+JI97yHYeJxfjjEQvC
U1roH0H81S04MXSoEWVhfUCP7RwaznJ/EQcJZj2fRA+PCka+FTu8vo+qDYgd1qNKbc5ocidYG+Zl
m8mDT3FEw39+uQfUUEs43SBURhD66Upr7BehgWRE8GhJsDMsyP2Do4K0x7IWinBPmEjm3SGMiNEC
ZTmKYUn46PmPbJlgSDDyMD6GNQ95HP5QleqBt3615uIYDkvmywq5Hn0axZ7qSpXYziNN8kzADxtT
OSJByGh8GhGjSKUNLTHAHcsOV2o7urLZnYs/gev4I/uTRFZw3RfPrEG+c6MB61Z8gJN1C7IAam6K
SxDsN/EOhMwfGVZgUIWbFg60evJt25WcGFS4istyyC3vA52/7n7idIVMz3NdGxn5fBdSBcBPR2BG
2YzlKjOP/NDr0q03YaQhrPcQ4fBvgnPJuR+LuXH+zAp3l7j2yAbkxu2EaqnkgtS2FOcNiUwpejwa
CBupqFOEnGbj2FzPTo6QAIod4CUs79y6NiYgEd1EpotpG+D1PIBdKt6OHlNNBu7Ey6+Iu5eAIg88
q8DfRRtbVSWlB290iSkFIXAYD8BL0lOUKmb7QTDVa6NlXqLtA9c08sLKafnLL8/01yskWCuWJrgB
pKVDoeyUbds5kF9CQRloVv9iHvuPp7tX3BfGhVDzkVlkivNvnpIaUSjxxSu1Sn1NBLRo3XgC0id2
9YcEWDp2fP9D0aBDLhv9MuaR0S6xsyopQtI20PsfuK2pXdbzDc+BDLoWfCeCyWdv2XUwm/ilAYHZ
Si76vlWdR7geCH64iZiamte2+EZC/Gzs2W4+aa4KCSserk21CCVK5ugCapFJ/UNy4H2R1xPBfvR2
j/ost0Vv2/vnQV7RxBlNZRw0YtRpdO2Rk3IqbMBoXRMp+LMzCax9La63mr+L4aMoBGYsy49DbywI
vkapdwvRlQ7DcOs9kOSL7bDx6Gdy6ESMZ3onem3ws2v0JkOJXJ5sUB5HluPaiiIbHCnSzjikrSy8
lJEmYAH+okG/RGFCo/o5KRwq/j24Jz5MJOOmie5E9ligsDhWgZckEuO0d3MAg5yYe1vobxUIv/2O
j9XQhQfT49nQrWcxCLJ3RUaXm4IdBjnLW9I/ylROyiFVd2hUBLzhkBR6RHqXHK0Vh+31cjXw2+Gw
V+t2LTe2KaW6umb0ErX4MdaPzToOOGb2g/cgKyvQJ4XidUiQ/7EHpxJ1yL0HxuA06AVLPSV+nR2y
QwcHDozJCoQzU5txg2nTvIs/YIZecoIh2fKpwkZ5zWa5kADy78WxCsI5TBFSHr2oZVaFoLE6Skln
ac82MMUKdwawVvpB45fmnkd1muPEKCnlMtMsjcnY2JfBp7fCEzGFvY/GHmSvByMp16Odp5T0KABN
bMA1VF6jetnnc0W1djDolOA5L0MCD27cgU+7XKKI3lo4xCBd4yfTzabbhLyFrZrP8yXZ0x4dy+Lw
8ICaHO/clHkwehfvXwQJPBEVzrXXYiHY7R0ik6Pjsc5DW3ojqysXNKQ5844PDigiVH2mmOHkjhIQ
P6OxVSrJPowwVjeZulKxtrJrBpux9sJgG5aBmvA7T/S3WmmEPCQYCSAHzA6NRm5NrIY5lEPdfwMt
+l1O4vIks1Z8M0t8SkT2PqordvWZUinLbuM0Cw5G5N+oyg2k2Jw323nm3J1nRelKkB/m8raDO6wt
BJoHtL/LLPxy9bUlqlsNAUoKdzzTGnGuUzelw6Qs2XumeMd1E/O8bErDgWpJtEr6CGVsB/bBtz89
cVkNXQpHiJC3yBfcxpUfLsggZOsPIjanRH+e2PfjWNOPskvJ0TCmRmoA7r/Ywefdjp6hwX6ocb9G
Dh/mtpS+wEHVvg0Llf3UClp/TjcTJxe8c8qtmseLIsOrKo1E0+NLFkjNtGexCafgLBEXZxYaFeK/
2ailgTReIg0X6+kjNINoZB/gK8k0QibYKx6zuToszEBstKh/e1cNVR7Ccl+ZC7MxIi1OsqAKyarh
DLW/LDBvSZFdIQ1q7KPoasILXNxidxs99aEZe6g34bnSvZveh4wrusQQQzvqkJIfs8a4bb5vOOku
mVsTD3LnsAzHsXXS/1GUZoBDfMjO+mipy/aTWUS5G/gQvPagVFLoDO2OuDy3hZCNmRplILOLwvDO
VGAvqrBGQY9k/vmGM53Mi1DxvoKsKNW10bh4P1Ekar7fhLoI45Rt1Kodnng8fA2Upp/UP66C9y4o
DOe+Uf3AgfScQjd2A70lfGjh+eR/bO49oEFDXpNuZDh2TUtSdr4n7MuuybMQOcvUYY0Nf/HQ+HSv
FgjEktGPtn+elht59ij9+PLtM7KQcXW3Zbo1jVnhfjifsGcC1+BhhAx89ifopaSQQaJyGLt8odUW
06CSXeDefYkOOjIoiD+9pjHpY7frTjr/YzK4pdXcb/FG1fZ4zz/BYC/8vhVveKS91ERplaJjYmvK
VOBnS4+GbCdaoGeJ/wVfz6xxC8SZd46T46l9j/zIgODPTl7D//OEihDmz95EzFpWUNoXPqTy440B
Y8tB6pTQLp2fghkCwoHX3334ykhAdaZ9wXqGq1Q7S7iWuiCZnZg2DM8QPvyyuqUbUdm4PLSVdKro
H3TfYY1U9uAnQ/bMoIwqBsCJqRPkDrLTJ6pNyjuWYq/3REdg48lSUAVaATUelzQmin5UsMH1G/fB
5iEjxCRY0ZFDVWGLMaNevqEX0OGXcTHTaD7SGnXZ43yVlcxn2HZ+WA+uT6+IVse51H6+rDEMBKNc
uyuX2AZxQ1XXnMdyTpvMiCerZiEyZVSkmxT43AAPbBL9rTG+IGjevSfHJdf8stbHcUhF2JomtEtS
0MgRQ8IOI9l+laAITNTczPxGo+5h6qn5OKbtUZq9E5QUUzwlIZp8cN9GJp0FYn/Wyd8I05SmSdXi
jw0ArzmiFUlwIeBFVlJ0nOTbWID4BBcO//29Ju2NciYAFE0puXl7ZXFtsni7lXom9SHokjPTWNeB
yI9XT0lJggSO1oD1+VvR/tKLmEXu8rQCt2XL/tIm47NGJ6ZZq5BD9n09X6l0xshKXHfBKLpEvlL2
E1o2FVEzhBJ4KVUli0h5/iDTQp2kSgv5uhmhiNQwsnZiGAPC6vEvg89UYEXXhf9GDziP1oWqPQWk
mfrsct91JBIbjpVt93zM36vEEuN4NgPQUXJCp0rY0iBavZTpuPID+U2+bYJZs8sgOrTaI/6UHLC4
cCConVkY17JVa67705rgwZFQxcGnRu0vk82x1OfovjqYesf62keCOgqG3q/NaMHjw4vMBUn0qjwx
IPXbXIK+826s3snhM8SgMhtWJ8+yM0EAeP2c7+d0Txn+4ZyE6FakN/WbDRH98/4eNJe7zL8cfX5D
/T38JalUsDujnBsDO1n/y+ctnuSLMr6iW7S0qOVWrcCORPZ8gdOSif7AK+8vsqmGURB8yOigLhOo
HqfHBWhMjFf+H6eaW87d/ohDn2nqdedOlzcnnQCmKS1ufFUKOhQ4vq2cSIgQVgGcoxKWUDqrKU9M
aWgx2SN1amfmUOywG0hheFEdrvokPNOp6Yay37qKAL1zdur9aq/2NWWmLLHeKg4l2jB4hAyJsg41
pgKtUIxVt4/MAiMzTC9OZqnGN5uiMZpIWTCXlgcTbAbba1CbwpkGNVd2x2k+O+rIe1rfN9cptBte
rDD5olIUeXdhp/z+D6zje6C0IQmWibtDZaJYVrqGotG/qZnt6wirb3VxykCBdljIu1FJeV0h4yfE
YWbja8TkgwVutrxs8QiUzyCL+rT470bpZB8klmAGSWyTyhYjR1fqJryh1iSs5PvJ9YAEoy9vJmcN
Vz+8UWiijSSY0Jr8qVzRc0V8FRR9EAhe2nbV/qJd0Eg4HpJUARNgZDO2IT2oKAhRba3nxAIjz0Dk
5F4FszKBf8jm4HyGNxt2m2qffB5jv8AHYzyjJ7u7M2TVgDMBkRjJpnSCTi2weHKLZxnQA4JI3Ecn
v5l3wJdQP+/iU62G2uEdIfBnnLLySbqqhA8Wzhr6oQfVKHpOdBfP6NWdUezkmS9/QgvigiifVowZ
v+KSHGR/A/QzUmQJiYG2sDZASyoC0TZ/Ve7hSYbdAoVdL/K/6CUvF6hX3FvIufpxrPkDJtsTYDa9
PRUD9PkUOSDK7hH4wi9hRFIDwg4qwT0d6C/pttSO2YVNCGvhpmemu7XcsS+pTRLS2+SxBtrbd2DS
z9yzeIaVvSnxhoHb8how22OmjIpRvE3qZ6bZh0cVCizbhTNA07WL2zGZUg5rGrJYBf1r1GokTtAi
Fl3ZYjr0h9JhVTaPjTGvZhy3rqMIASJuGWJB8RC46Ut69BVLczcDCs57LHXGqEK/bv2Ru9nEWwBU
Qk2UuDRpCMfjSxPnoGBaOoH4mXE7to0QcgNQeryskAq0p2a6pqQPY8BduJr2oFaxd0/3vUvaCBqe
aMvVdCOrSpOymgbXqArhoNBXreYvnhus/UnDiGlA4ieuDERX7aP/1dsQ6htHsid101CpWYJpRSz6
BkBKEx1Q6adHzxuDY3wO4IHPWkb0AqGHLErn7Flxn4ysFJ+aRQ1BxyleoocDiKAfBJmXOLHrLjH5
uRbBrj1CL7SJ0pgewLHyQGCHfVwxoIZMsKmgVz8lrTm48JLSzxP4CrYap1+boGsRdz/IejaNksG5
LpS8Q0IAdj/wKvNUBM558HNZvw+cIocDLnT1Rii3GoRMy1kCaAjpshhj4O9sM1TEwCl4cuiWUaIL
7ZupTFsieZ9fYu5tSB4KVfYUasZBD6BSM8vzYrO8YXQi/dJZYisUt5BgfACSbm1z7jFDk+kPNSV/
FcFBwn+/R4mpTGnrunyoh7+zxy/+DurMf8SCiBCJafdxF+oGl409xclUlDZLBczxG4tHw5rjq8q7
ezBbCt2zL98LSpcYQPjhsSABoqVn5OWpZOFIAMm+UBaTNAiobYP6QuWIylXO1VjXgWjNMP5Lgm6a
k/oOmH1GQ0ARa0HUNBzfNSTdN6ldN3V8z6W6HbCQCTyuYpbML3+vcQNGljKNykICo3t8SRo2FnwU
3eSIrAXh6014VqFBaMelUIy7Z6ie3zqwKtr3EO4O4gVbFjlATIsZY28IC1FD39MoK9qqjqJB4ssU
SW6DS53JlclnhrPV/2yerPmdoEItfkjOnSgJhms7qJNOePjZ2WIhPLzQ8jU7G+W4yFY4uhD0pGer
AA0FumhLQNp21nnUEZ+rlbw5b2ri9g9NpuZj8C89TdiqcLdetaRVy2NWOeNzquTdKwtTNjFZogIr
aaL/B+5T9EhHQrkngAf99UsbbFdmOOrEIj+Ykec5S/KtrDPX/c2A8qyBgX7zToIa3zWRfHVaKGnU
T3H9vTLViBw7USCvA8mZpuMIcnk4tFEEO3xG4xdsaW2wu9w7A5JMLLCOs9Ew8S1N2kbJqRNM+0q5
tbsSafDi7l87XQovBg8S8EAAqB5fNjgvSW5+ude3l4bHhreZZDYsa5YdFdCGwV3CQPXv7fKKO+h/
eABBJYCIzxda9uzokiCf/lSth/jOGew3GWFuCjBOvydOtgQMJ3jsDM3gSqnwxnzQGjoXKprQ/Gyx
s5r0XDgNrUdIakVveH0ZvoUQGOzm12y72sXXjwo10RROE2OT1DbGf7d38iFnxQT04olVc1XYad2i
nOHCxAPUUU4tQb8XbKuRJinPIyQ/oGdb13vBGMlAuRp5nRWYby15p8H798fpwuHmnx0xNv9AElv5
uymLgUBVhg0QCEjdsTkL/70qe9WLBywgfQZ7RJd1oKq8hQbh0Yfw8c26Avcs0fVXo3d4AsKYR9iv
nEdBwpc0fUdjibz7fclMXNd7DMDWDRyRw4PwlQ2cyFY/kN1nEAe+0/ZjZ148xBM+GCvI+8iUnIP1
GH17XO5GrwI+c4O3mHaEmu1mzy8cvDY2RKgHm8D7gldR512z02XMZQ4APwEzcmbv1RdywL1GQIAd
pxNcsVEdno6MrAqA09sI6rCvcYXBi9LZiJcOSY8T9YOBhE3+DwV8rt9lSxbYMJ/yGqqQ1O2aNuuI
s5DPxW8Fqihni79p+uNIRkryd7UnjHGhRTuF2dSzE9+sOLSrkZ3nTunmYNPBpJWx4d6vOmsfExJU
SUAy0IdLeoJ3KXlOoW7WUPgxNuWLkAt9jkL+Yd3DIF7178CD0ITtlh8GZplVMKqleWSTtuXJkgiW
iXxF62haK+npJDE6mjeLw+FC4t7mid11uul5lIZBDO7PVfwhwfR6qYQq/+Sx9kTdhEyaoGf6/pTj
v6veO0q6Jsey+0pfG2QHDV7uxLS3ESTuDPdFIRKmW4k0ZfIpFSdaw9RcOoVqltIGUYNgruGo6CSt
afIx8Sd6zXA8ymE5334CXTbYW6Uv9Hv+NCaDzxahUwpj2cnvpy8v8fPcCriEEuAUp6w+1itdDJ0U
OE+Nsmt/yPlxFDLII7i2JjzEdWTe4+xC6aUZKC3n1oVbeeuj9eIjZiXomQRxmqllljvgBqBKctdH
/KRM0ojbYTjY5kXJ0Ac8oMHHA2Ah6bWaTpOlsVPecVJxO4XDI/FYQbCi2oGOCY8uB6zeoubaNrNr
kLlp4uGqvyN7F9Ho3iK3hIpXdJfRaAAcGsvKB+Q42NT/hHnFk0v7X7a5FNcnLpcPrJtWUySwLaZq
8BEV4AuzEQllGy/trByDlwU4dT9Wb6TvXELqVZBc9sRoT3/vDNTuSS1jc5QBZ28I9cuYH6V+suly
iDozc6FWAuXFvU0OozlTemb6iI5NCqk+vRvI3WAx0AWf99CxtiL2oVodJaBw0ZETRzr4uHgSS+vj
bGSMDPhv9EUgiOmtRufXj6moWehYuZiTJFXNn6uybTRdUDqWVV5FfSWSXTYBEAAiW4e4szBRKmhI
m5OlC366EOkPxgxBmwIObuSFEcZ0U8qyw+S8YDUr9ryfyIlDCMPnTYhgScUfk310ouByGKWQmWlR
VgeqBj1vUOucBONo4nNyO1S+OAU3becv4AcomSN4uafy3YwsnxxWgrzOpSI+ucq9K+LujGdeQQV6
2bBn/UTOwEl6Xq9YZL4lChZeUL+vfeUB3Huy2zsO/ep60ND1EWpMJtlwgO0w1JZ/Czupwq/wg9/p
04qmfUUNXgi3e4EYKR71dHW3bRzqpcjOh5X+dmOWGprmwFRHZ+Y3OJZy19NNc31ICsuOrMyclbCW
0l3dON+zvRJURyMIUlcwLZDqMIrsFyZI/CcgHdZ3YeyWXNneuMNAolOnyh68TqXNL4REvcOwSyZz
DlP9+Jx0YhMP9YTshlC0g2ycTrnze8Sd4NlWLy1f1wPAyvhIKgrs148ZDS1AYeKWcFvAvixYJGQZ
FUgzJtFYa428RQ7+POHtsd6ab43ow6yi+ZO+f6NjM/Ef8DbrCgd6PnLlAVNLVwa4zyCosbCah1HP
zAMxqYhsH/Zsc3olCoVzwJM9ekj/gPh+In5NMwhK9eQ5DMklXysmrBJRp7jGCK/xbgNiHYP4/K9b
EylsE27WFx4VtUResRyUBfn/UuDxqWw8hxBL9nSC4UJ7t1Qh4FP5Siz6/g7xAV4DymeQuTf3L0L2
5j+n2yBWFglXQzDzvv0nRr0OO7Crb8jycDgTWZV/L5neiJoU3zJdJNmPg8CexzjMq5IZT2fjArbM
AXhAQ+gfEwOjwsFQzGEgLWPiUSYFEd1mamxzVUuxSRHDVShJfaWkFWDk5d1WWyb9UUHs2du4SZV2
U5iooZBYFklFiKO2C1PG7LoyYZksFGgBYNGPHHSClF9egEbFUS+xX/BJ6cRU8LUoKVZhaI+LvFfh
ChrzeOOnHHild5MOGkeE+eI9XVi3f3PVvxEVkABfowGpcmKSdHr6Pi8L6niISwschEON2BDYNoX2
8nDT7eBadbDvfAb+OsE6SqlyU9yR7pO5w3dY2tp4FnwCHeUJkr8ZyuA15S/g/Jx3OouWFGLt51tF
N7tw+oGENZha3lati6yMd8KcVoCmCpWfeHb4SRMfrXDdFbwzSCIaMs7hCDYOAcU0n+6OAOtsNhHw
Mm//+TeuPnWxh9uimGWc521wUbCw1mYlTvYM/GazYXq2QWPBkyS1Ypam1TyhQf3Yn/2Nm0ym1o26
+upBSr7ue3PNI1/Orh3+wKAzgxZ5uJvbGU+6WQJjdYU+HbgptJFrcZn8wpK65KRqR/aZj82aiAR/
/5LuEtgL/YZd6su+7vIGIFtAS86bCPaW5jU8Q55RQum2Qq6Xf3WPY++QJ4B5YPlF0CTKId2tzy74
+8V6oXjkeZf9cL/FS92bpnBCwktShVcvhhB8Yxw+8ZfHZ/bj0TNog9iSf+3dJgOanQ9k3thh2x6y
9bqPAS/0E1lsp70S8PQcFgWN8ysdmb+2nKmZoLxeAk1nUygdtfubsXlxdNhuLEKex9sBTbXCLuSx
8ts3kZQJPSLQxGlabSlKvuWR2mr/BH37yxBtRQdq2r55TNUACpyy87ytYpanGSsWHlmhv6qNDXWy
fgLlgXUhDRMhH3bi8ls/X2zDjNhy3XJiddZPYTrG89F8WrY4rJFRgsJcu4dSXZvvksiW9zsZOsjW
qRHCjvRACE7OsFM5/WeZjkIBd3dnaCSfeyzG5AiURMxtiCMhIjicgR6YKxK6Ae1tdK5nxfiEo5zB
rXouxVRtsedLWfXPKU42pl+QU1/3D0V3D+6bReFFIUW65RJp98KSx8XXAr51SwCarwJgRCx8014k
JdA69l/Ps8kR5/T7kpc479YbHep7BKQrJUu2KRN9+xDoe5fth7kf01iaMl9pX0NEfMKo+rTXUJLB
6MimsgvuK+Tq41ms0V2VcfN4snwQjsuYrxY2wvGWS00DE/7liYbM0ol3Ap+oLgV6vqV4ibiyb909
1Nz2NFpZcEaltMs/r58ho07GKIOOn1dto/mLyDCyfKKYcNoePqP7YrHPDYAxRWJtIYVEujwq6EV1
WTjf6RJvEPTGxBTP2Y1Bj0h8OxiVuhZJGsyPiGe0XIHD/N8x9TWelH+CGLIdKFPqTy2FRhf9sgln
v3bDdM194nzyId4wWAWqSjACVDcBi+Ti8eU22jPg4krifiqhS3vcnkdUHQfw90gt+D2WQNfV3AK7
qyR7o9CLp2dXyvfLjQ/oE2r4lnmMLP31X1qMYjdehRbcLQUyZE+Q0u+GhMz7OIco2S1PvgBwRG2W
Mep7kqYwy0X3AhgWpQuK7JS4Kh5HdzQhPVeJdqR5xS7KULetFoxAXnNP/b5b6dDgTVd7qk9s9Na4
jiXz3w6Zhm2ESCoZuCnF5RVdBn4cYhwfNppKd7uNWImx5ghOOkdCOkIBkxTTVip/9IoFiNJlhqLB
pyj4s//vpAVQ1vVDGvFN98d7QrDpFmkCfGbgXjsCoCHAIqe8wu8aU6Ih6K3uBBMsKbDf74dDJmk/
gg/iYBZ1q9Z+kmJbGWBlwduRri2D5oetAQ/fUSnz7atkUAXILNniAp2Gda4ot4CvD/KHzJRB6tGm
82kifM2SraWP+1EHDs/4yTsJLavF9s5v4PTZGkCNSXwp3hQF8wJf1cXykhEQmErxDL87CYoElmyM
3/5YCpeHamIZ+ekI8bONLjeK0yuzrX3rVPyfv1xH//oJiIFbeB45eFEifxCkbAwhyc/nwTDMGEST
+ryP6dnA2JTziKfg4qxGRlbGDRz72w+9qen8cdzzNCIYYnw0iRrKhKuZyxkNRvgB2bb1rDjBsozH
LwzO/tMnAExvYfVlH7k8CyeEtGK2ID+SAXYdL5pFj6Tigiz7xEMUwEtibMfm9JtNz4nvEeiTUJBu
WoXMCUotooFGji+grhP2P/3y7xq28ms3GrSdBhrmKT4NXCm4cFpORYrKAZNxYapQHmRBKCj92kBP
Ywc5bpU6hAKuOWe02B+9p8HtnFYX/RhkLEo5zBQkJwg99ftrFPqn5MVuuFeaLyEWI+2Kv9Cw6eRn
b0QtoUvXTKSEeXKkUmkqLDWgWJPsMfXI+Fm76m5WRZn9/FLoA+N3WElOZBPWLCGHHIGADNdiQelK
RUxpaw0WyyNohLQfKjSMSBhuA5H4GT6w0p8vMXtxjarzEgnqkusgpj+WRANjamPdKGWiz9Q0MBde
6j6i+5DDi1sO2QqpPA6COAdujVIeu2THXK83AgtqVW2bD8q5xpXDxAZtGMDXaCCRMCScf2s3f41s
4q8/PSvRbQX/bcM9F8ZwpVuJLuIEWu15+1o1MggmunrM9Uwe5xH4tX/Y786XBhaMS1PK0v6eUNkC
h24+qJwKXqC56FovAjf+QGkUDURG0D8d2D9FEvAp5FMEpOEP/M6lXXZja+F75b7gniM3Gv8zv8hp
DZ8EAs2HgvzHxrPgcFPJOT34FCCn4XJeITAiHb+qTsz+vYc/VPGU4sb+BCqx6pYEyxWNt0jxP4Gj
oc6AuyMk+NmPWyfP5nIpmmSSMqI9Y6I0PDl8JnGkt0uXT7rgHbBgOof0o6Umqn7z6lqw+6qZCdlZ
dvCL8JTRMRPiC8DfzP7oEWodS6cvL4g5VHT43COQvpZ2ysvLAmRJzvA6URIuicaqTPMcY4GnmrD4
ZxBaNt/4bJs9pYDSTS/ASleK2g2gGjy2QHEYGGepJlwzCZKJ2KE3Yuq89sjcwTbmdnXZMCgMMqmM
44CduuliKfxgPATyhkBZbJ8IIMLJ9W5nM8I5vfr5cGsgGGTMJ3L7VwCwEU5nBlUkuiFZX9OyFloW
rzoAZj85mv+a6T9Kh6t/VfQw2r23+EYUwx9Y+qjoNxXBXm9lFMiTlAuHvzcBgsNyNLIETm0hMBQr
aBTu86W2YvFJDfPRF40Y5RSxmvWMLhZi3GHsNiCDU790sCB4vAjOJzX3IzyZU5G/soKABxYkBTdD
+YEcuhLrthrCL7OygFnEvAZOOSRo3E2jFgw7NpHVv7PhvHqCTQX3OxvJFI1s1f795jzcpZyMvOWZ
T+jRqX0990WDL+ZwKYgl0/RONxi4gQGpO9cwUX9YmleV6wMrRV0SXWnPlU1D+XwNZi5pRcMlhmQ6
+PtogtvAXbh97oRhH5xlbKfy4j+xM+YJeeZz57U2IkVWW9jBberloTGZ290Vm2QUTHbzDpiW1vBO
hRT1PnSk/Ye13qq/tkKf9b3uY00abtYmXmlbqaWU5zYm+qKcnTQZ1x7WRKDhJBhv+ncReOqrhtCn
Y1QJhjvgenhxvtxl2KOvEVsg8DVB1vThfpl5MH0NgQON0bp5ilZniFOpJfcdR/PqVShxqEGY6t7x
i5pClwrehrApsRxnL16loTiyKEqaiCIUupm0I2Kc6FASLtRQbdMMpkYBBRFQMDNwsSoKpcUC0oTd
HRZWg14+hCz+Ul4mqAnjhn0q/5v5klj9RrvfH6db7nkshNioDmnJjDne6xGWfpMW9ooNedbEtT9F
c/DydDSLg/BjrRouKS1CswMqJ2u53HlyXr0jBkz0X66hvatmXe3Cjd4ANUAt5gyrcI9sCPw57Xb1
+coOxeupsBcCmRd3AuqVA/jeGgFm1uricR7/zN0p+Vo9SXYdaCam+zG4JN/i7qfX+GlUPQnk/dEv
3crlGU1kurHcIkJn5Xyho9xDKFLbG5yanb2ISJDysFw1llcN924ySG4JkewAoz35QSWXLTarDLIh
AdANmxD8by8bWH1Hp+EHKRsZBML+960SBgc1jldsgAw169PViTYdkx45NcUhNmS/nNPPheIHjU6R
aiHlbNVrDvqXcTIXs3H/eJD3JuOnUznCknNlB2X10vJWNDD2c/VigH28QVI72OGAu25mn/N71VhD
/AQIueLgd3eIUrRl0QWG+zUa0wsW7R98nUx1uYL9OOf6i9RL8kInANTjRH+ZUx0E9VGG5JJar7B4
grI8hofs+BqCxk077SYKmgAGd1h+DtN2+juZ24tl+CseW/lfYYUHayhx9NeLuon7XgQmiDI/8Sno
HBHMn1wB8L3LQ5BtvYZltsUzvW/zIgNSp9npR7GueZTMnsN0CUajnA6oc/vxzsj7Pfi4kDlo9n77
x2fl1mZi93hNqK7lxdiap3FqeKeWWp0Tqi9TRhP+BYR35ql0+nOVVnmqLUv/suOPIEw5Btd0Pqnt
57dDn6s/EpssqN3OJnL1BkbhwccB0IJ6YIpvuTpYsItZZq+o7XmUeh53AHF9cAlIXWMtGcc97Hi2
tMtToJLkqnvW1xvFrO3dFK+HRZPNUEltdo5v3dDj27DQCxYSaQthxyJnSy76y/h3aafeOaBibzS7
eCcSNGGgqAMgtKCU8UvkqZnIuw5PXboWmCvT5ripsPo20n1NX3T4zroyKRrBZAxVKiWu+Grstr1t
IGi3RbtGtJB9EHOjd3opgejT5FXtcQl7sdSlSmKw+DWATXTQs0mYCvtj1Midd3GX0SEiGXiRkhIe
b57NLjn9OosrZ9sqcUNrFdOU4CbsezJ/Eeg8fU/E9KRLhVE3Ctn1g9YKUiN3EA40019FEO4KPIyK
IEjnupnKj7mKXkkEQC6lCpbwD9krePNO26+YYGgMgoayqi+UZ5cd83Vs7kgOKCGMKbuFMn9Tg1bf
MKUwxVH/5MJVCMnbqwdA8qBmZYBG+j2uTojKCNqH6CwzU4T9hiIBOm0n1vRfdtFYvX+77bSwl1Bt
AuNcSbg8Al/1PkQt9IpwYidO6Gd/UQSEFyaQKB7slRouToEdd+QfbPyUZqKUrPSCqUFdV1OVhCJR
Qf8GDVPXTYEsOZIOXhJbJOWh3Q2hKqgy7ls1pr4uW+ss7vJvfToBsXwe/ZWlxt1tVM58sofTwfEJ
0XFxl4vnYEij3I9gDKWcECTdqBXzTbBg79LVErGcnEZK6CHR3klgPiKvLxPqdQl4R8c1q9pU3OnK
jbMjIHQ0PaVQxCQWssWhSAx+IFsik9qN3ZfXWwkcqEfSDQ1wlQbtFhI+Q2OIAOPlriOVR/6n8klu
8YcjGQo8VlOO0ZXPdhL2D4nri0PXlmQb6fO+KHWoTm0lkI9VeyDguaWRVnrSQ0sKtL0OoNQ/pNaL
wO3WS1fchdSYm2u4i6b5Pu9S+WazTwqtOs8fNDbdm/QfC97UJOltMdwIolqdb9O7kO/ysKZiAYjj
SgZrAtiggZtn1IYgr9X9dxpPU54FgUMFl15hmk4kywErMYYvQ3Uu/SmE98aCgwBx2+klSs+2NOkn
fo4+QRSG/2s2VEGYy2zMfXYBhUZ3AJY82OmlwGWjuyu97arckoT9Nk+J5JZA2j2fq7amHTIhZbnz
I/bCsPlNwiOo5qoGJNQiTdvCPAdk/azIuxpA35TP21tVjTxJmiGMGZOvr6FG7gSqSr2G6KlAykpI
Ns91m7185qFGf7jTHmTfF6kRogSkZeob4m50GFXM2jiLjmeOjFTLjYpTMOK2RJMB55N6+DbgpGbo
L7HYnXI9Sv9LEqCvIwmbrwkagcuKO92mSE6LtUnIL5bkooOpqyOMgW2ai/vkQjqlc7qK5yoYRRDO
zTlzL1hTLTzezPCrq0YETslzgaKB8smKRznNlcm13awl6f+z1K+frHw9QUR8B+pkQPMms8YBXIzH
NhN/QLLsWrD6/E5ucAqrb/1VSwaaxzUKa1brq7ryn8C1Sphqfuhfz/CkzpfqDIg8wBAeqb33SLzk
L6axH0RaP02fvSc9XxMVMzKL673yrd4ZDGMtD36bC9DKpW4u0JsNrovHjIc7HGOF9/mGWh2k0QDF
5xcjLkymEikf+dY5z3Uj3h9TEdb4o+A6uGuRf4CQaXARJvnYgMv35sRAMjepwwxy6VVT0jyAEEY+
oryqZVEob0+x8Sk04y25sSd2fpAQ0fcGjCHCUpCSfbRBY2Nl3LW94JV5XdoPpsWBXGa1SCWjn7M3
96LQNju1MVGgFUOnWCfWkCr0Ipcz6MJFlzsxstxTJ+O3CStrEO/tUoV44Lw+cKh2D+MzJI5IXbE1
KGLfXTfPgNy/VRufLkKgMYlaGgvxY/76eaNq5GRjfSA5p4SOl6pxtvUZ1Z/KfNhKudm3rmdOCsU4
EOa5TcVPi+Nrc1OiqPDXLWtd3SNlSkY+wCxSygB8FRWfNOwwWvYnzEoP7P40aQcT8MgUrAD7iqM9
PjX00+tQVw1pwFc3YbJZWE57Zj8eooEOhrlOarN315ybLm4QBR+onM1e3nfLaTJ2kKz7K9kSWEtc
SkfKrv5LM7F7nNRd9Se2r8SRR+imWJtJJcr5JNwKLaeNrKQe4b00MqSRg1H2G5tnlWqKKA+TU9iv
b1vcCc4fTPfKoQE4/ZxbkrmfZijIz188pKScX+xegtxulTLEEgkj9JSs4NpI+SbbdqFR6A7wDEww
dg41A6HA1skQ0HIQ0RJo+88dNLQSmLxaBPsfzBczvKW1tNSlGLNrGEDZk5GfX+TpWNv/uyk7cAfw
iuwQP8Syv2VxFYGBLOTkB03bl6aGcj6wcpAEFOD4nOi44emyq20nEuACcaXnqEiMpaBQatEK8lyG
W49NvfJqcg7EjDlbN/yVRnA190wrd176fJTapRSSY3osEayFd5xm7G0iirLImuSVnwg49yvArw+f
bfYDc99ndWaR/i5550Q2uTZMKH4HWlE41yIqZw40uLSfUNjizKdmV4ShlhHBJ16OXtMCXLkQ7GS4
hXm6uUumUQ3wvJU2dZOf9CvBZJXVoBaWS5OE/u5x+IZZfCaA73AreZtkB7dZuMp+rLESX5wdWTvN
gHQLeDXcAznnxq/FeX2RAXAWBi8Nil9EteoSPZBwjNrZ1AY9R1yJe4VIJ8bvUaGay98T2ldycZxp
hbwTDiyaxT+EUag/FLCjZwfuhrQqgmjwihClBPWrRKNwZe0uIZ8RIIAdhQxHk1UpJPzeGVpkwh70
FlwZ4VQ5W2jdtMLFOpzibE+GSMimbobsx1y0dMmmWkXgV94mL7++NBAqbqZ+1nm3b+A1XTxW6qU5
DjmA7jGW9woKxCbmMQ6ed8Vy7/KjjTAbqDjXYadvjIhDxWyq4wszPQc+z0PoQ8tytljnz4sUbhZ2
Lz1ZQ4VzzkaHD/4SLZvzldasSJehBYK0zzuixB13LU2dx9VLlJ4o37J0cbBFh8lSlG+/zIPO+88G
GDp54uZBooB75jgcT45xOmz0og3moFJqu4z/JS0d/gi/PU5KVgVjWTe28eNLXcJR2DYoY3QysfCi
yZDz57L1sYbqtwR6KVVfgp8VgF8mrO6dY6SDW6Yp/TESqWQVSV+xlnMIX+optaazsqK3gzMU81ON
boU01vtSZJovuROI7X1dxqW/K1lf8ojnpbBtffevcoLuROj3/4BpXJoEmYqaXv0PE1FA6AGcPXGW
VOxB6LlYpPxRTqxdholVNo8N8IN7pyFi/zkGvLG5HIOFfzce1BXmp0yy05KuUyls+IFhRktBrbq2
HWQnWlldQ4AMkQkWNjPTOmEQ58OTMG+md+xD6oLsI6MpE4yJCAus9mI1LKF5qZ7xM2JSslK28INZ
SGQbiJLLedygEytqBt4RHkUlDFWt7pmGQ/Hwb/OPEzaCf4ZeYxtmsj0Nluv6iTVMsxwi5gbomgBn
KxwrekOF5CCi2WQmMk2m6PyF5vjpMOJevq2p8IxobkEypnvHPrlOjVytGwhHEEt54kbHm7ZsB4SY
h2oGAwnwzxpy+pq9ByFBG94gunpurUO8H6Lz0oB0ii7sIhoDfveJAm5YHtxZO8FVvQZc7hvpIfq0
XQT2RFQ5oPppXLL4prfu9twmcUoEr/RH/8VR8GSZwXrb3ZxafLYIwIKJ6EvOELkP5NOE2fyaS+eb
mZFgMIw+snDNIzlpAOJv/RCdKtuC6Uf315tGvg30RXJgqs3c5G1sbyb/9RtVjq/clw/avBtlKX9N
yPVXxs+7ZEcbLisn5KZNYKD2c82NObupw5Y9MXBQe8OO82TWT1LXlrOUHFhs+cR6nCqxD2siSip6
1BCVoMW6FzQlu+lTtl1OF7paFiQif3sWbun5ma2XrEKbcTBNzy0Lfh53GzKZBxCYg302sTeE4aYX
SfId2ot4rNT1BMw8xfCzxlgenBoBOx2A748jYOcExuASvfjc+WPhyxhVFJbs2zNlLrLMBYoG4b5y
/GtaFCDFNqTatVzEemIK3ZKW3LoT/GXS+FkfeBz8PvdJ7jc3srZCLHY6rlg/Cjm82Q/QJKhntvXL
MjU+0uy+7vcOQKo6NcVXPlKPtrD5bK/0G4dqk5mU9pkNWk+tE29YG0hJdK6ah7K7UcMO50qWE2av
a3vn8uDOLJg0fUQYfCTipZYlluODkIFa7hQXyjz7ctSeR275RSOmRGauqmlxAIJDtHTvNhkc3sgZ
dC5PKW/zPA94HekhHzQoamcDvN0QIxbnUeVIHKKFnxaHGZX2EFcOreu4lVmV/8OdQkm40WY6hVuu
rwuALTxKuFuwu9L59KmE97vtutsBqfR1yySFwEttjU+fWjTvnH4/CStw2IIFpCjXbfEiF99jy3Vq
qrjcwFU3OqLl/BRUVgNvnU97+fnRfqTt8u1mbWO7JJbKP9tqt30o3sR9PSFwZ+cIIt4YE1aWMgdU
XyeIjwcJlp9wA+uvb+OhjqwI1w+lcLXfhjU30Y8+3g1udtvYXb6LfMqOb4hUWhYCRcSobTPUZGrQ
sIdmUigRRhPtZlicNPqOnsIu3boHK8p5InY279EeCbqti5xD8OSGfBJE3qGFTYahzUyM8Lz6hGmM
rL1ipt3Hadoif2DlmU+Y47ED1wv6zXT6QlHle+Qq6v7+JaecqyX8CTKwaCOO3ULRpbeGUJ30FgPG
O2sG72mmh91qBfNJMUWLdcDlncilrt2P0IxdVPjXGvHAI2QXhepiC0a8o+6pXfDYUyEdv2KH6UuX
UNdsmr24GbhZ7SZYAfnZ14FO652SfdpvLg0vvf2CmxSHF3JTiDPCZYwxPMhjRn7h9wkQX4fNZ1bB
0SQpYD/e7c5P9pK8mkh/sLTEg4vssnayFxO+xrdZf2eGmpwmlr+sKljlUB1caN+Pe2LIkm8/4V+2
8ffwGh5QVsuN232u2cTBY682IEtjoFSkOYxw960peoGGgeo/kP97Dnl8MDMMPPGwQliTcb/5Yn9b
bs3WRiOeIkLzQP6zFF2IFaVW8uN5Uqp0ejK2Kynj18fjA7VIJ+/xtONyvdZSlooitNWaJ+xkmDxw
OO0CLoBH37hcvkpvFib6pz3/3TLqhiG9lZKm2juRBdZ4bAohEoB6LJ+HAA6W3n5GgNBTSugxzczu
nDntCXAL7ABeaCK3dzYeJY6klmuw9Y93SUXipdn0p4wg6asgjbG1KPCV5a0fs5dvPp85RJW1M52e
WGw2TQflzCsFUDvvT23/FE51FdLrB/+TNEdbbu91AyF1EzeITxNrJJ8KrDO1T+ZHtlQNVzoCdUZC
W0ub+6dws7JlOqpQcP5U/h4QNVrBl/l53OB+Rxvr0eZoH9azeCbW47GGpBghxsNzv3SotV/iKFoT
WfJlfPFIN2TTWA/pioqPIuCfoX7/jttYW6ThYJaPrbflXj+To1MFKqiAJA5S86MUjgkG9Knk8tvS
jGE8loTc1zat1B25+m5mqmOhzsJch9bMk1wLt5XOudEKVt+wv9RJ9GEGvoIN52qDmXzuxVdSY/8U
kBzLV9xg4qu84yY6uLN3r1cnM2U4ZB8OKKHRy5nwgqEKBj+amnNH4zoKC5Uzi1ZKRwL3jBolJ4OK
KuQ+liNLZdOV3JiSE7RR7ebENCZP5mMglers8spXcncsQWXwdSgwM2S4I4P7p2nHmjFoc97uzpz6
tgKLwZjsUVkfQKBK13oLiuV8R+sqdNk6pheWluOgaoep9TXzJfIEEgUy6lU/TBnnvdRtBE7VP59T
rnrlXcEAPXXgykX6hahsOdna8of4ZrjQyLJ8+xZOV21kVFWYBl9dX3Kk8XEmZ4wS0ZGH5DWwsXU6
cS7Yc9aQ/pcNy+gkLo2t4qi6vqREHixXxLHKz4Gc7iHATkgLYabDy9u0J0TplCgJk6imoxJQgHLm
hb7aXy7779eYCgDmte5pL9bx3/3KGWhK6tTcX3WfuzzMH3QD8uZL5WLXvRWEHYHhjqLwxpA573/Q
iA+9ofwc27BgxReCW9gkofdsD4Thyvrlp+Puw15h29llv41C1tMMPg7vSnhOyiL+hkaXs7KGkZ4a
eVNoN0NQjG7Mc3PLFXezeyqvPtF+NaZQhErMIKxGp66vTjdZUZZNmJNDUvvYgQn928bieX5oOJbT
A6r/nLzJPoZcIJRvBQaCo0zZr6IuwHID9S4MURAnm57MGjL3BYT28MgIKNTjbMvuZqx/2hHHExbH
1cELKfz0PAkHiP+U3FYegXlgSTHTWSrifAUt3BZowFoFbWMwI5+fmQmWUw/V/kc+tgjLqz0lxCWW
bP9sKrm8Vkz7ty4vN3RWqW83T+zw/5dvtC8tHVL9u12Edd1hawxmdby47sBLrUsflvEonZCLjwLG
noVOUSUmnHYLYR1O7uMKPfFBZDGJkEDyeKySUcrxqlpWs45M/G4FUhzo/2pw52+MlOMbOlIE5fk7
ROrOTLENXtwgg292oD+xSUgIxvb214P8VqPbPAy+lvZB9Kox7cpLQM1iRej9oGfT8sVuCtNRfBSh
qeh9bBqRvIzYyDKLkeOBQQ9qoXrBPDAlA0CCH68XIIM5UrN1ufefxFoUZoveT2Am8MFu3+V11yup
KQvp6Q56Oj63Ah8iYiGdTz6cDhq2xxbVwwATH11+mVesodWKiQzc+m/B0PpH5ty4Us4vUYnWEVUE
50aW7gpqfEYYAHjIQTVE2d739e/Dq8wkmMiiOp/9hhzwtIZH6RW+YmDdwhyYbRXdOeH7Lsm1Ml4e
uRVyyYFOF4d72LX0mXU7K14EyfTCT51Qs4wjwrutkZ9fNe6/whdMWGcY5K60Fi984I21aJfeb2ZD
cr3gPTIpZD0vsC5O3VixNQI014Zx0uXFYB6VH58vyWBxamXNNqGa36XBJGG33l5j8yZJqVqpGIvu
Dk7cWjfvAHwYMAZd+jvB4fNF/FD7ds0yc25X4mQF7VuwJXJ5VtnXkgrdPzV6Z+UixosU4Fg4/bu0
OANZyNa3KICLMUrYne0P74CqaR4jfLXmDr1WFNbO3pd6ZSrPBFtFnF8q9RuEIl2B6Ce8H2SMX7O/
oNtV54V/l7vHqdSkpeGAW6TLmq7xJhX/avpyfZDLMdNO4YVHl7Juq/EYTFET43yJ80cQQp8ROeF/
nKAWQecyejUOPkkq3LhIpwemVhqvHXPRNPzC+tqgI2Vxrz2XjET+/WNoEOZkvTwFRmIDMpLByQsV
1QylZpLHQa+gTkj2rDIGGoQA0BjCoZOLTtPMqTRSuzKeXHVyjeCb1XyQqQrhxuG3asgoQ/u57FeM
YU8cEdtDKurri0wIC8No4Gfon9VoQhyZNS8XXD1jKtLT0goyGq4ev+8l+imw+Lib524F96S24+Fr
B4Hpb8/S+XAkmrL7BeNNiUBqzUrX0zeUSzjerOeyMBWcvw+MaCx9owtoxccLbB0HUJnw2HjxRtV8
a6i4JSGROc0r+rA9BAwrceqA5bw7xf2+uAGIgznIbprXqVDXFEubJEfVJnvtrQyY1WBZ/YpimDHC
YhoUr9Tb8zS9QKuT0GfHMMTEeY4UzK8fTkxwQ/3CiewlbxwZkCQxKPdweAp9OTx10bgQEXu3fEs5
by5ac6wTVP0e72sGH4ek3kLoiUmWNKF0FPLDN7luN7mNXa5/vXHH8hUgS2Y+QbA5HYhyfWWR6dPA
/6DDoNer60V/592ruEQlwTwMs/e2zDhzlsAcx5x/O75OIh/HCDZC0yhRs5aSKk6i2znYQ5bNHNrs
tcisua7DWMCZcnOUMchnwRgESG8riucCDHbT3TgGknAMssGVpVceyDd2+E1819wVf/kH9ISKvky7
6M+oYsazORs3VM064r5Q+SlkJhSmOAufauxkTuTqIx1KiMScvfrNr+FLCqshzZUhqi49fFnB/dYc
w1a3RRs29m+3hQ//aEVdijmIQnG4IbroTLqIBfi9Q/ks2JXDfUA1GMqmJNQiou2DkqwPCl2Lp/Ca
FYPa2CsHVFl9cDPJWcNaKjQjQ7OzVzlYYwQvRzV1n7dmWBLhj/LH2hHU9VasS361o6nVyFtuj13h
lBqTR9yRsMfX4krLQCPTx6JUkwdywTsVBmPIUIgoQtyDRvGYN+3owrDpT4mGE+HUpXlw/6mD4h9P
BPSuxuyh+7xWE8+0zxuX6cJ/rTgaac9v0T1v921j7t2axmjX5JZTtIIC0gin0Mr9ejT2wZwwgNSs
PHwbV4GI5ctdbnaue6TfWOcdPMiNrWuCuTLNSuZCgGiqapHXKArIl/nlKinwyq2bNWJcxVaSH+Ui
SZvusAgwSAbRY2ud79sFLl6CQ+zF4xjSaKtk6SAnjWLhx+ktm0K/q1FYWbNJMWMZQJ/ArZqPWDW7
YR3qAl+PV09skMTpWdC3QQ8Z3KTJyl429GAsJJKdDCq2EGvvcTp6Esn67lYZeUjdPPM0mWCs73Kk
HPmm3i5fSGOuPR7wQDAls9k91HpsZtp6NwtbZCGlW7LJDdcEA7LoBCzSikyzLBD+HYj2H5aRP2iU
jbXrfZY5VQaYZc8mCzIMWkwiDrHp0NH6T64dRxc8/SBOuaxlpgnuTKIdGrBVC8CmjNKGkS/muC3X
v9/5qb1CipjjnVna2nXDW/TATb3Lhxl0lzjm1s+PkBCGPvN3G79AlJtNkmF/TOy1GsgLhrcmevbh
6OLYqAujGArtJ2AkPyLH7fQ0qej5j17L0svVI75m20X9GkDkM6mQKUkCeUmM0aT1UkrMqz5ZrfAW
GvXEmAY4+Ff2j2uICtMvD6uBv+RGbe2daSpuvrXO7aE7wTgi4rzeLlYPIr62jkwilcP90zhTSrTU
37pHB4XaEul4dZcuW7pdHozGvONRhwJQYFmqklaiZlfVTHmO/aRV3FLXW8gH+5zesJ659nz9WOZT
viPX499Uz5EybQ+TrXxdSR6D/ui7dUZe2cXbKfkasIe727tNp28W3A6Ppiv7FQEK82xnouI6EUOh
74qiX9nUcSWUezYU+GVHooELYTD+J0zbw01Pc91F1VZxy4GUCtlk6eGwoPL+HONXLVi3DnmLxMMr
RA3VCYAVHVEdjB4kFjsph5e2LXhnWe3aTw5BhQN9eEZdD1rHtk/YPC11R6WY9vR76aDcxNJ1cMHZ
11bOFmvXBxBd2GUnki4XF8Og+DYiUc39DMWFTr4pJ7rq+6jIY2MEYhpfyQ2qSse0ut39ghlbo+ct
jGFDo/yiYIqB3j46mIws0oD/Sk/dQEkcpthsjsxhvqUgT/7VDQitADSBGGBYxcnbTStegIC/ItGs
QjvQN2ahiFWs4F94mMI1yAEjEZcrAUots7rtNC6eIGPdNqfEPvgtb7bY/wGXfU4UoX9mwWdSp1ed
MFEb03JK72r32fB55YIrXDf1ALoYXkrBkZp1ZRxBMJyRBUSXC+Htl141hNYKCW8IIJBiO/S/Y4sx
sySmtdP4b4GH5nZXz3VNrZ9q9/1BWSIF58RAGPu0Ctl6kxfJJIntIxaG2NVl5R2rLD1qZAXBaPyQ
SH/nXJZnQqntoCJPstd7D6gCL5vzsEUT2krM6rHv5V2WVYs8jgGLv5IWmyc7lsFAnaLkZLcjeMFV
ru5B3ExoU6SeNMkGoMN9ZyiTtveYqzohtJtXsQkA/pZPrTI/UsPmjeBn5bgTgeBht0pmwTzELwNC
rI/lYDe7CFOVFAs9uM4AJMTOyCUG8/qayBqV9m+WYTCr8an1HfS217QHnJmBpVbyRJG0kChlHivS
UVP0zN/Jl1KTV7mY2WsYwvB0hNZnxO+BhmxjxXrTj/L8vm5kPUeUfplGM1vuyeOZxrDbWICdvKBG
sJqdmq4azqQHhlGWojYkIJ4OL8vgWL3B+LeUsyAAmDEXAsEjeXnY8jcfhL1pLqOorDq7tIM6UyHx
3hAaL719mzNHZ2yT3rUox8cC/gkOJybZ4Ky7UK7ridmeWcrVAhRG+eEx8M/EwdwdDqdIGkYrPYq0
Dcra9/9SWv+vHetaS5+wDYZR3tja8tA/mvMjWksT2ZsbltNyV9WBGMQmkmSDMtMFsadG7Nc1SVDp
jGE4CPXBFIbdqVZh5OmoUiCGS7Y1VajuEUGOfILB82I72N/yZ+eoSesVbLtvcNsLO2WkSMZGaawo
XU7wY3m4Ift7Tp5x9RnZPh2Y2orzyOtFZNBiSNNquQTYV/tIFNslmYZ5vkquHVBlEcnC4OvO30f3
Wkaw3+Fw2Ld2W209sDcgzD9SHx0UhIeK/qGBWUGrG66vQqmdnX9WI/PZtmES9X8usj59PvLOumAY
SbOccFQ21a0Uou2Y9ifkVBxfh1aJ9p5tzknYKdQfacOTovwPPWdm0MHf2x6Mx99ihX+NYzOFVuUl
TJTHVkbz9CEQlSVNy7h+T7vMfhW+DQgC2E09qcXd0VfngQUedUExXFiETpYEqNP13HkP4/QXBaos
oaEb3vs2wyIFKFKC6uYKQzNafvKhjQC58H2r9I2Yw7eWpxK9REuG08pZTTaIx56VwQQ1wgvwc4S3
Li+7mI3y3d7j+NACJr6ZE9Sl+OC++MgDiL3KUpHHofNcGx8LqSJ6sRVCekhl72B2ehdQp9i+ao0W
Faz3hqbR6BvRL6CJPVvM6JlQn7l3qWSgnQSSFksT38ssNlxDfcWtSMXX6O0ki1R0fhMAPR2wGUzB
1O57DKcxKjbLwbVxpcj4ORJsQm2B1ulcOregRluWd3eK7aBfw5Pu/sUzbfjDk8jy9sV4FIEuRkiq
d0NwAwav0F1BDYNUuOrgN/8s1Mp09c21hWOG0W3aSyj1ji+uBBk9QDlEcwj8Y+j75VKuhchAyCZX
9gAOZwkREh+oEcWxY2fs14lW4F0aLAYsGbPHQOE5mneC1zor1f0Tye7zhQgs+KvJukbN1i1dJJAz
Qpv1+04Nb8eY0AUMgPvHQElkm7jQdCX4TcoXztPuhdLJdyHGxuBiS/Lk8fiQ6NaOMn41dj/dTkE+
hJA1p9oUK/nNvXJFky01a0aICTz7aAlhnxTUeaxyKpkz+hqjEJT2N6YF8skfyN08A4SSSNKiez19
yexLCIoCOjykuI2mO5XrXbhR92oolTpWGp2AhUr6AJcE4z2+5Lc5qDy3LUsim0F8ReepJCc3FKay
ZmmcnoznKnwAP7jch5jvNWnW4LTK1mkPia3mpJ5ysAfFKv8p17nVGOh0OazrveM9eIb7gpW10nf0
1J/1hpH1hFexp1ALd3sU0+vT0OKJfbHemfLNKf/tG2FB9WudUPtl75DiMSFo8ME34h8ESsUn69/8
uqf5N0U1Egr/BPeR1NxqUP7dEr9KdDZS0hkA7XweBJ9qrz0GvlLpN3BW7EbtKNNLrs8ilYvRFY//
aKkfaJSRB0CGLKoqD8bkwsYjlp8sUoj6cpdFaEsDsHaOz74XNHM4FEdW+RoI0FOd4Qgj0GaAyre+
7px1EVxCBS/1ApN6pgqABxy1QDv0WhLhjRwIhTnAXUyRc4OhThTAjmcprLNxpRfF7nvEYWypI2lg
p00ed4frDjzyIEEgfCguv2HmVIdY0hyr+hFQ2fHxg4y5iFrtM9Y+twUocCCK518UFxoXRGYO4R82
MeahDr7MNaRzNS0acV1kIIzPA2pkrHauwkHBf9uLp9O2Y6O3oo4KjA20lvVfaH2ponrDksWwmG+B
tXHgSUviT8OYScuS5SpfysvQdBlPmKiaMzgJuQVTIDOegWw/6mK6OKqaoCWlkO64MailUGN9Hny3
HqFnv8j4jqSrZ4+jP5nzoYVdcbV+fkHvdwR7WAklpaV1xrmoEv2bTyqNv+emyhG1VxL+qWZTHOj8
3Z7Mp47vzChJiwWBJTHm3zi0xLNCFnYFeY6NOs/CayvBoztEqigdCfszImkpGsaKEr7rZXRqnnq0
xj6u+aQtkOHliCAgrdbbGdxxmiMVshjIok1fO0rdjjyA1+cD9qxZirAKUlwHB7dzQyBxNhqsPmjy
rcA3h5GveV3Tdd/Vi3vAJu53naveiyV4e4BjOSEBlFJ24uqNynwEWRdwn4rRmYQsbaBTCQsS5yH8
yD3jLHCVNCBE9reFLzD2BXkcoxC4YdgREzA6H24U2Mni/droaF+TXVft8JVAEHykI5tqTGLLQqNt
5z/az+AESp1n8kD4Mbh8oeH4qcZPUVZ17hLUIeJf5Z+D6eSEgV8pF5GYCwbux3QDUY9eap7ibo9d
6r6n0XD7HbWpd0xWQCAFy6QTkeZ8h5tU1PioDEg/kzgKQYKtXHe/RAoVnDIZEv9d1u1RNyqDL8ZQ
lUaFV9aMbgrJQWnuUuw2u7xeB/25MNR3D8iq0uihWf9KSjRWcloFMEhJ2ISM9dPXF3eAuMTxO9Ks
RS1tO28fXB/IYl6Zv3vfu0OLSKO3PmkIv32saExVPCXNpnWT/86RQvtIJI0U/6iLlLDkL1EtmLII
wz9CP+80UMQw+9BuB6sIPWRK68DMjGTDS2B97NVTZxrB9dNnNO7BvKs2WeGqHscS2sKi1O7RNITl
cy51UutquAjqBV/0SRqFHtxEpFxO9qrvCdnvr+0ltDWxLqyO7YLiGyoFxPL1qE15gXGxoC8GtsN3
bN6j97lWSkU3KeNctWo/diAS4Ogf3LTzTDU+iWgOb2ISIeX8IKloIhRDYXTlZbFEAT0R08ZQ7VX1
LnU8kqSk6+FLth0mvM6AhiaitXB6rSwJO9yQQ06CP3pGDvLC/XSHng/ZAyXEKbrXSemS8pjitZdC
u+z82KqALAM73TzKAfpQpXroL4fZsiMjbVp08fXpemmID2N8s1z80vavYZ2Dmy6O8s4GGaRX1hDv
d4uC2J/RBfEGL7Zp0RtJNEhkblBl5oEyjRq/HzWUlOLd/WiW0z17wLGZ6FJHigPK+Isbb0G3W9Hp
aoHd0NFzMEb7fiDgGLIxyExUKQGQkxkiivMPEPP6tmLKNbUE41JF72rS2GCNl79MERFe5WgHBp+R
gIt+OfPaLWlx5UNgcUBJw65z0g2ixrNidlS3Tb431hTzkhmNze127nBhpInSPIUwv0FVOb0MYg/w
9J2osgWN19lnayBZeKMO5MrpgBMkkBr49xFbXq70znJbyNwHepsHl8KbnQw+p3XsYDVsRX71zAU0
ZN+clBfj+VgRwmRtjjFKqHDVN7COlypPxWCsapdu/xbvNPa+JuIVVijEPLHkgZhaQOBbglCYPAzE
huebjL8onmDVna5AccFK+Q6J499hPzqSqQ0CvkTbPdDiIYTEjoMwjKUGW1/LKqOPnJbdSBSppGYk
/rddSEdJ9l12aOxi7VbyVZE/Uqw/eZcVfLSdjjstJpOpMsQNOpEsxINTIwp2PBfqk9+4xqCoAeGF
lZjxGGz0FGOstJwHl0rNxKNWLVXfNqnOCZoh3gje5XUZRp7d3ShYUeIkDS5R5wt703veX644grAi
++l8PCKQ4DzA9W9L3fOOrt2J43JNNidmzBwU0JvlrEM0tIzClR4EoFDwCmM7hcyDEFuP8/D3nNfk
wMmLSII+c8KzZDWS2TNXjsxOGhtv1j9yqzWtkv8IBihGQLFUu+tnZjuaIegdpimenXAEuh2zzsYX
kWPfe0fS2CXf1jP5vFcsabcc7R4/ltvWyZEpBNtyEIefjByvZ3tcXywPGfg3YS7y1B7Jnk5VNjx9
50KptAOHcVzkk9i5FZDjznjabeP23izYKOFVH5SQBqdl+f89pj9vSbxKcff+vjWSZzjNQ7gLi06R
JgBNtpAUyIOWXROounftmPK53KqYk1ZxS0Y3tp4KQYZpOI/brPiNJELAQN3a6qyOb1t41a2HUJ07
3q0VUA9zBad6+I+uw9b9q9L3UaiTUl6lB/ZjCF7/mB+S2EvkQEU0DEBNdPJrIpxlbA9ZejP4O+S3
uz9bwWdg5xbDGC2NAa/ubG69f0qZadPyD7G7tN24+lKppAG8Y95/NHEPnHrzcrSbatFOuauMPLTi
vvvGUIuOFBzJQbTiKGHJvkM/8VjqFt47PSNAFyO+4aALKczObi2d+WFZDKM2ILYC9wdbWNOw2mJ4
OmxOgmdVoc17odxRnHJKaK2zATPb2Ug4k9qkFK6/izxoclyE/zggLXEgS+sEpR4Q1p1LKmjrjtzA
hf8eAjckol0vLCzbzlo8FlbgDO8mF266QYat8juxp4uGRi13yXcYC5NE7aoSnsioR2eM1MLfkBYW
e9DHmSzZLJ1opCD5XPW0ELFGqpAfxQdLZn98JSR50gCvB4wYiBkZgKOWo44+JORES3r4IC0JsWqg
c3UmL/6KWVIMkS71LEvbLE4Fvf2cx+307QG0CQUb/U/lAzUIVpO/fGgMLBY3CgZ7z1EIXwF/slZT
wBbt0MS2KzNYKByDKwmcQRI/YjfBYrsMLe3vT9Fe3dP9GuV6WkFHubLIhMT59zzh93+/0792dGrO
R8rWt3F0Vnhl0dGdK34dXltEAf8zPX37myR3GBEOY5fQYrIUxorHlPYVsNRgf1E1yfOlwVYxDoEq
jvjZfDVcf2pfrydSs4NRstir88P8qf1HHq8/wqiRJzYRNV3syQ/P2V+WLNnJIzk22Cg9DDs3q3LW
26Ydn5JmNhjwrxVNUQXNnTF2AnVvlz+lAH1mjyjEz5K7s9zvNnCmvnJiXgY9Q9DXos4SAycJlPED
eABBXbk2NGdhU9ODmQkmfmbFHaclObx//f0uXN+EibUIwVeRpt0zQd7onf4L+gzBIRXOmVebyjAB
iznYHHisYpRDJMdIgGihB5GeuCNh7Hmgwj8uIkPMPDmsFwIiNOmguECUVocNwjrJUk3HijN0ZTEg
Vim3Or0lvgzLARlae9B+uSd69BlBSMRSGGtWZsVBESLuCrsMbu11W2yF7pZ+vVU2dDx2+NE4MdRC
CZfm0K8HD/sX3M4YrEPNU5ktxIVjTAhzlEFB7pr/vda6jYmLC+7MEmFD7/ftobQ9m53MdBiAC9qg
BaG8x+bR0qHeOnKu3voykhEkdiSwObcGiQHfzl97r1UAmuuQuaj5R0isuqF+zGWEXE4f73cIw7oY
4Xp5X7nh/Y3ZsPzSOXgniR3avAvfgSQQu5O3N4k4xp0zgpd+0OW7+VwjOzhp2xfHVWZCh+mHpz0Q
XYpzK0emP72F7uI8Zx5OnG7oiF98f1X3dNrFTxEvjmlrkytUUS5lQfQevnlwTHMxVroTnj9czCwu
cTgdsIt9WgX5RH2kYcL/VVYmcowGuAqNXFXjk3yJr8YqdblrFhgmEhLbWu5Str0lysP8HR7n2Fe2
LuAUEuMkRS2wrPsabJHgsk3M1GXAbEkLxD7Lw7GqU7347WntbIGMkB9jHD3mjSIYpHpbHKJNb66g
diP9saPpiq0+Agpjgx8qjeD7G4TQKDKHxBg8NRKo/idNTInau59E9mBkvv1xY3HKKzT/VzvsipHa
9XstwYULQPe1Dm8wUniPAE5EZRr9wyoMJZR7bNC/+NcchdK+6nK7BpvHxHY/tdiX0mW0KWGGGgT7
pOqv2A0NCjTc+uMGi2znIcpcbWGAdEV0tljgF78Yp76rnWAoqQIaVLu43EkaCv7KFEbCdUFvo7Ur
RuL74E3HUAuyZVVYwev1FsPY2SiS/uV/xU+6B6FJC6U3DrjVNZcc6YBT/LDCsFwzWEw+SClFIwe5
6l7VwnHh9DFduuNODKRnyoVZxsV1Zh13czujA2Aaz9647+/x4tT1+dtfAjHf4wi8dKcDUuubAVer
fKSe96xoG+5dCx4pPnxuo5sHbNAO9NSp+bpdj4QROJMMsizNMQHLhZrJO0R9iR5wqrSSrbEB3TEe
slIC2iQ5WQ4v4Phb/6d1tjO5nQhZQ+sMZ/AGH51v7zPujhf1dihVfxWPGYNMxZVOavLxP3GixfM9
+TRmE3FfOu9NiI48LXYnfQzccLblp54MXFG0skCPD5Al9QC4EQv1GOcK7nCSICu22tCYapE7Iusg
mnYg1ZSSD1HhONraJJyI0xeWzm6u5afaw0R9Oq3lZ9fsYBMwJLolxleg+Mxu+vbWT95WgU96dNyH
zxpEJc2EDD8k3V0+dTuYfBDQwZnY6IC4mryamlNwmzwdj/qURc195UdcWoCDCJ+Jb43pwZtgqnvj
wAHCbVcJCfcY9Z0pkqVHtJaDYzTHKbu8sozxkXRe3nDglaSos6ioHO8ZZQwJ9n8Dl74T3udvDA9k
LqVH8P3XMV4oOqwPTFydH4d4U5jZsNeGcD10tgJypLzMfUjn1vg1XmoZkUH2GrLG25+OzNa4TYOg
1+9ymOYxMvjd5zvR/7oXefKCmgM8pCMEo+nVosrthliEnSd3fCdwWEHHcItpi68G4KryxEpJyDiX
iGuLFb+bZu2XLBi7oGBetwq3dKx1B5iznsnpfz21dXDtkQqyZjWL82xq2EVIV9cpQWQ/DzBEGx1m
VTHsUA4PCK/RplIWV+GicOWwUJbYAdiqTU4lDmZzOjh0nAciQr2C6seH1DntBIg2DQ5eh64Q2PbD
aYMiezC9X9e1WWcouHlQFG1oXcvuT+0N4e55XoMDOWZM0sOOVIkb9/IuQbWa0akozAfNQbehIz9X
FHxq6ZVTFh8Xst47spHfs4L+yHjWBMN7IeT/bnX8PoGcZMsnzuT/R1N6Wui8u/uiyvsPn/vEjhIa
9L6jQfzPA11TdpInGqAbkkg7743+FGPvdo3rDzJVqlTZGYLZV+SKyjjmheGbAKGKKHq+9aBMqD0z
l2VCDvjSVlJbGACcO1hfrVVSO0PABcz4W4WOsiiNQwqBKOv0g0/JWFkXmkBb2i2Didx+D5yjTSmh
cT2ieurBrWQ97AubmM3o63sIjEcLk2Kox8jZYyeemgJSEI4Y8esVzt9DSNpHCKXBX8bHsh//XO0A
0/bDJa6wBH/ipD48CUDFzYRwz7oZxlZOojSl+sx7LwBHBKMtiV486jb3wMqZy6IBNESuxckaqzJj
i8KQg4gDHUH7CtkJ/j5h5iZfUkhwNqrrqYClxBzFbLCT+5eg9aVYH3l4ZboqLd5w0kvzMQ5xDTdw
duAagD2rAeh/JSVuBZpEogQTUxXG+XIWqu0plm/tjNfMhfSHKAHuDJNUq8+KWYWqGIewrz4tJZl7
X22MVXaVxPK2WhyC/udlfIa7uVoWeijsgtvJxk5la4A6qatugbNHk1KZ1nQsC9/LIaSuQUKnCAT1
YPnNsTlSRbI7YJlnYC2IQ4/zygOQ8zBwhsxNJyWZRKzdg11+Pzjdto3gdGL3yitwSJcjFwXe77xP
16U3bAH1/dQXhf26cwfuGmKQhrGQAqCAb/AUPGr/5GgXkEknIweAZjpkfbUAmpMSM5ER8MguH5mW
RTHcHMxgp/0hz0Njqgy6DRzvMoQwUWMp+gc5FI0CYxbUrglf2+vHklq+TXU5D6LDRobe4fw/ijrn
IDRvP9ZrwfoIUGhHOMCSTt2CjWgm3wdAGSBcxBV27V+ZRUB0RDmwj8Nsayuc1auZfKZKr0pEtcsj
P1otIsS5xm8pkUvCNhwK69tkxDKvCtOB3MLq1NqgFULlkWHtHuTpXXTgzgN/s3wfDc9JFahB2Di6
Dh3QxKf8huQofJJqAQgNrZzRG9uqgiD9oyTCD03mI5ghVwrayc1cwSA7w7U8amCd/wLKnKgEmYao
jyiTzsAgC3BZAb++Pupc7lM2SiwrwRVUd3thCo+J+5P590nfihaSzsqigS4yGH8z3otZUOzdRmxH
L0fPK0aW7hJmnogHf7cnzUvMKmU/oWJiQxxQFXKyqPhpaFvtX94Ccow6Nzf6HqGNGZLFEv+xSgpK
yRmHuv9s8nfbAXk6LbJqxwC8X0ij9vtHWny1C+ic5t7bzzDuMDG2Quau0lF/KQ52aXD/6beQRZo2
jE/Rk54QlqxQk2NRoSt1yVxjx5Z/4DhvlIYOdLPskvkcd5hrZ2YBFSwuCiB3Ltkr4+Q5mkTX1E41
i8PlDguhQ7M9gG62PCZ/6c2CxchYG1ArGdHzWq0DYU+utdbo248auN3dwt3zPycHh6B/sn4Dys2p
zMnGlQw+wgPWWnb1STFWWpfQfe8oIDKwjiiWmoE7m9XTqq7x6A5WLADkYRLFxrpLO5gTSCJcYXvI
K+8kdoE7VQlYIYYd6cL8/InDeI1QJUiq8HtOK4BsObgdJDB+wqbA+KzXeZnLbDEjZeRni9ZQCHgj
5Qq3F7N22qPJAAMXg2Lfj/SCXBPVyqF22tsJre4LM8LVAyZFFWCRgVQovywwrou0n5i/87XvRtN2
RORR3H5l//fAz99YkMJ5FsDT7wRax8R8caVtb9vjkhJBzMtQ4BJ/TQP25RdBh5iLznQcCUJ6Lxic
00tKDLtirUbxuIl0DCCkjxGmkUQUcztviavS4HHZ27IMrNHYhC3T003RwayW5c/IILhQT8vxyYdS
EPW+gtk2I4gqBhduDPhQ+IfoMcR+c35HsUtCiLzjk+43iu4UmrRcqS5xE43imjp7Kysn7Af1NxaJ
iI8XdYW2CjTXieqSeEHzN8sbsQKJNc0doj38YefAi0+PVJTY5MtcZVy/RcMe0et4JR/2ORqBK7uA
X3ZZk/DwNXlpODfZ5zvv4l1gEbkiA71qdFWK6ZSbIIpWsXRqIw9K9gqKS+qxOR8IyfsTsD2j5O60
PwIEUPX/fTqDsaC4CZ21k51x9swmF5YxHrETE2LS57aOueZ/w4NIm4X+IYaQ+OmJzAXk0eE1kwEb
WkFp+SY7chsZIxVLfByZqN6xUAlStQglycHZbHnJQjahTNZJface7ZijvsRbgLK3jq1n1aRSl3Vg
0u4CjRh1puaT4eTo5OuWcQoDbydByPqVzrRjvagJfLvzf1ZzYx7vJPeSL7BEQgtxBFrCHU/OPl7r
PMsDpezZigx7btrtOjw7qYJ4Gy6NAL1xjOcVDjvrnjZqgsCwHNHspsZbzxC6NJJGH0qeGUbsGE36
fhJwm6Exkjuda2IKJhSVi9IYYEXfcjoMfyqR9jS0OxZJP770XSeGCPMDqOZvc0EYQ8jwT6RKh048
Rf1EpEZYYwrxkKUJaiochU4O8dTDExvfepDFQg0UVY/pcRRKQULe80fC03oLsBzfYOVTQrnMfMGf
4FpdL5nODkN/UNUBwqMOs2xDRH+D5mlZIcbJrm3+RT+9UcfeaKXPEbmOs/2NBb1ejCCDWwK54+g1
IOmvMN13i870Y52z1lDno2F3fdT6bB8CRgyzSBUZ2fMjbRDwUD87DxD033p9AJVYH5793EthfHzL
e7j2RCGmLu+jTq1+AN5ObFxgqM/Hy3cRGXuTnQ4r61RkN06/EypKqrAn9Ao5foXYfq/7jeCkcwzf
cqaieNescOrmVscM2Kf7TIRtCIj/vBeDP7nm828j/qIHHMPftIMknx4bsdyYujttoASDFnJvqFGV
57y1d38mGq/cT6UnjiAVXphYh/KMPuVLHAnC6MiEbYEv89//LICTqnO5t2K0VEjNTCYO//Wocx0o
0Ome7zUrmc9HElw4FceyL4uFCYw23FwiNnSus5dEBDEuqyrm72g92438vE+UqiT0hgp36HQP1ZGE
Xki/dv9xW2/GeT1DyD3kZMlIO8mEBwp5yVISN7iREz5n04RosA3Ilh08sypJqfoZBVSER1RSLVQc
2Zb8D0sQyjGTf57aAEHmonFcDTb1OsjqF9YnRqRihFmZFxUjgFHX6RnwJ9l0BiFfkzPeoyIeyGGy
sputbABH9l241oQth6oVBZAb02ncMMzToCiRegx0JwjIvhBFVq7wUB4rQDRryDokPRLmUq9H4pud
GvV5LA+uY6RumJt7OIOQaWPAHzVg3cAAujaTeaZd5Kw4UScrLXD/QVEGwlC4mENachuQgEZIy/Vh
nd+wAf6uImM9ECGxMxag1yiP/iOzbLxPuc7LequArbIDdwHr+6djxNaH4QJ8dpeEtxU86Bro/OOt
uFBVhpipqS2bsaD1mf3kN9WIwRHYHrFq9x0c62TIEpLW+dSMEmhBENEsXy7LVWyIfw2vJTFGj61F
wwSpO4OzsKQrJep6v1uCilCNG57bgAlSxT6V4Hzxcu5r0kcEmGZclsnprhIfLxYikmUzVCM/hGxt
lwaOjVeejwK7HFTjfx2PqfgAQVgT8fRCyNPvg63kkiR1Q2v7Z4Yp+boHBlzXIEnToOtWTWnpASvU
iFf59VhZX1f1wCNgYlHyYaLsrCEHryGNqlil9Su1knJrS6vEn9Bz8VAvfk94BgBSKSMkWBnSdaDI
YSvUtHrlXfH5n0HtqgOFumNjqaET6K/w8XONjW4NUORJ1TG6LTDcLTxP1jDM9gnd1ITupbsv93AH
hHR0PSG11NaUB+iGE0UYRUMnpgzC17Pdvf8bgvggTWwjXgCCAWEbMfL7VgdlKN+mAYJAaFliQeKX
Ej4SSvPfVyI9RlWDN9XkBJra4Wrkcm5KbeRh0fLbnEVfLvfRua9TzUb3GFyOe9NUBednG2luzVHJ
SSoBT/Tjg/9Zu3BdfoU7xXeLMiU5OyIb82tacrJddcDhu9e7fWkqHhMlF9mouSOaBpgOxDq/Quu2
rL130XHyy0hILctmZ4wATTLZ794/okIiWWFM3RyoJfngC/t/9ri5989GjStEwbmTTEj+32v2n+O2
D9HumVKt/htHfSHQoB6dwdcAxXpmdShko8aS3JQI9WfqgeIpp3Yy2AqHKu/xgBO2ud472NfX6PTG
ABc2gQDdj4WnqwSBtWfzQkZ4osL0PdegRtpDjsLcq6a9i1IP9OV6dbNTIMoBOaicSn0NR02z9Wxv
klBYDHvl13JNisRpmWIUBsha9XFYG5vuGjvCnCDwokEz1gdTKQZ5vPc++qBsUgjtGBwVSSDFgKBb
M6La1iKmUf7v7VULYCeuKaV3e2UebhCcag/QTdWf+R6aRsbHO9OwpQsPlJkmVl1U0LyZeI9RoXG+
VybM16p2dUh0JLAvQoRhMHHC+XJmu/uTj8DtdjLzASAT4A3n7MXaOucQTAZJ5VGt79vwpMBtkAXM
AmeU1xsGzOOGbc3uqi2RziZ2cZcpdyuLnb7GOBrddK0Iw9yA0G2PkpU+FlS5QAPaOsWt+hKnLrQw
mbtZuDUHvuehHwWgvOcX714omQ2pK9cqL6t/bwfDbYwqDeT82KbLtIoXqcG3k3IJlj11PeBfwpDa
ijl0cFAnxpSt3kkLixp7El5XTJLpFrT68ZQXSCYfVT+5WOlyJt9nMxK5xp5zdv7pHvCvcfY58DRG
XANbRBrZXfztG7r35JONFa2IJGPCl17o7OQ7mec7wpVR5vLabOZlygZsoXhKcsc7US1k9mqhoQ3P
h1LSJNlRfH2SWzMoc/216iW7L9OaeLZzSHw6hiuDgkyIxjE+27mfttmRMVtPPk0jR0lWNoYgiWXP
m5Sm8kE73uFjVUFnhUP4SwDrIZxt+uT/eXfan0F8KNZg04EcWHr/TVTZoSfUKBWB9vfn0g19IwxK
7AY1zW1CKj3C1HsyH9g1cfsNsOZfPq7uaHLRlUTP/1AwhKWyMwmGJWeGy3iqsvpd+wTS1s9GPq+1
CYgpQGP6d7lYo0BWMVh/BSvjDaz4k7kiq1zjL/9QtDZIr6WXP9lBh3E7Z8Vz8OJkPAnbkkMsMpyY
CKWyuLUZ8j+dd1DDi60+EwmMDYBnLQX9q+E5eY7VrwSFecT8/BlMSZ34/VWqE7Qq3TkJ/KG63M1G
1wEC+P4t8JsOvB41EEXuRJr1SkxJxbxSaBUWJLnRINsO58WV/Q6ly3qpPxTIELTglnUhLp03xn4R
aFz8vbK51iQU3OS3OBqw9VYmXdr3QMxSXIXwSPnRKoiEBv0ZCRT/CcCf8067vozQWApzGQfopOTL
udBO2HmobT5gZLp2pV3nyaoXr3ATQbZYutrCujx61sCB3hw0aJh5BrOYufwgZI53miBtB3wRiVZQ
7Q4XrAT19IuZc/T/EWmLKo6113dmrl5v+htcNfku/zXnohhjq4+6pGCRZmtB9yR3/20yxy7He2qh
4LNZwlYzWJt8Uu21ptykpuk+5pI67/hu6zTwgwjEE83yudjMylTuGN53EaUhRGqOEN/ckdjMW6f+
cz608W29qDKiLrPWozBCp7Pf5w6y+rDKDXiqloIC4P/NuP3X2upfqd0bxUWObu7UIKe88ggSun28
4t//090U0vPlzKVjgSpXW6XDXLJc2cWrm1kxFp3FnzPFBUT2+tBp6iyZbyNDovs2BJyHcwvGZwMY
514MHEmtMx4FMEN3M8T2vogRNNiqY3taBm9+zHdnWyhtZ6PjoPCt4SuWrg1Rr3axm1gk5bW1Mw9k
ciK0kWpQeuKXwCA3rgwXFM1A3DWOptdtAPJSeCzvp/GMwg2hxO8sVrVQKYAmXzQXJNAz5eAKkUk2
rbFAslEzQDpvaKmB/pl49sCGBxInhh1wsVPql0zytJTNNxJksu4unC1ItKzlZ4jpBGNqmacOS0jU
KAsSfZ8t1l4VuAkClTKOJlKN8+lswrk6PYOqFSKzQu3GImREUyJ6/j+dAARn2NMPn8Pduxot6B3U
IuAUeVMtm+A1KOSMA/uht70s7cAGTxES/tHQfLIXbekFojEnRkTsti1ysulZGaY9NOuEiGZd9g+W
nQD43xZcYbI4PA4RVTCUEQZSexKPpB1la10p33bVSJcTs0zK7aGj2vreZkHppMvLy1HH104GR3iQ
9b5/2JlxEMQsx94UqVm+oktpUxcDybigIu3GTT7QyUG62esomkkhCyY/uGsMbNh3y7fD8EBa4tKz
Hcf5wFtP4QAUmK3TzbPYeTti+p6M86bm9TGGj7O1sYIyqw+wGUpwTSJ1DjW3XRiJhassGX/ZpvYR
UTbu+9SjQ8jTV6P9BFwYeWD6vWAxJGH4h2llbvrem0/4P1IYDz7XSQeiZLPyT702tWDHze0T3ylF
yfHCIbMkukmwDeijaGx58OLIg3rhT2eHg0mxeyB41gsfvvt+In0sJweC7G3vC7rRy6+qMFtKsRu6
3LljGV2n3PNDwlywwsKT73AJvZ2Z/wd2Y7MtCYSC1EEP8KV0LlREFn8sjglA4dsb5ejFP5bPF3N3
zeyzVw4lPFuACa5nXRuVaiplNaWonEGg8vbLCXD2WPi5NlThubTNz54Rk4fmMTp0Gix0ff7Md68n
L5eHANyzSFwuGBjVicaSUsSFRbbjo03UDueQjsmAaLMv2PMBiLBLyAdSL43QojXql24/tOt+iAMY
DrT688nV5DUgIyRLJ0C3Y5NP4Uq8+pYfRnKvQIYBO8GHu+JuH0hVSkzZlazFiezGfJNLwTxTy6lr
OtJMom4NhYbXnEeaoUNIC1N5fkqSXBgjcxVjnnZkJTXPGsVsnDU3vLzI2cignq+QpK4irvZq6oEQ
PYQ2VAioA7aWffxVIDyDmJpytwGJ5v+5SS2+ADX7fKs73Z7pumxx/y4mWBvh0dpJb5PO4grNRXGa
DSaekrgyEN1+uYdy8+gifuGzNMT+RNpzG9/Dsk165rVBqzceAwQ40J/9t8ulSo8bfPx7SQEfJask
0CYohe6HoFPCa+8G56ZU6tqba9IGaULMeRxshpzi7Snc6aYUD5y5rBDcSVopYminN1ZBBHTt/W23
XJdHwRoatNcni0xWelljRyBgLKn7ElL4shZYXkxIQXGJBYL+RxXzPglzeEZHX1PjElpkibhfsHzT
m0hu1CJwuyG3ohd2ZgtCcKq/1P/NGTyzD4v04GUZiTCeeU3WhQhzDzbDC3N1WkmpFyUT77zHX1SD
2Pg2N++ibkHfV8hE1Wpt7TyPMOg8Tqp0Of8/eApQ/ZJcxTXIamsjLTiSStqY0iVER92Dq0nYzroL
NF0VsBnbiYtvUJUolMqvF/xLtCUXnLOtO2OS0MUt661f9NWcMFOhsgi40gnz0PGcXsEvEHGnIcxP
o8XGkWDnA7k3mSFY+IhFKXwsz5z1zTtD+LKPVsNKCedEwvRsv13IHqdjtIRntjSSEQn1os+Ly4Fr
AMhrB0kdekzjBauML179Swxq+V3tu7Yxs9ikSDIdJMaWx7prKnQgON+pZKm6lBsKoXmJ7dczvAuS
N3c9kV26SOtNDRirXx7JTGuauW610svlcgtuY0oHuwO/UB2xyCQCsYWpKQxRoawHIcQ0sK4ok7m0
IGO1ucSKEKd5+LiE1oxWmGCGt+5H4Ftc418H8Sg3Jhvp2A9fW+NaVf4Tbjc5k66+862C/4fwdcX7
HjR+449vaa74HhU6p0/wdPwCRgnIXAR2SZFVeSOhkHsxy0/TfB1CV459KhOAqeJHY6d/4fB3Ht7p
js+3n9VFSQ3eardoKFtlLWAsuYU2VadRmoGINBtoep3MTTHwi4yRZsmQsl+9QHJXfOQRdB2SLBe3
562kl4v7kc5GvhWNtdQDLpoWPprQnpKXdYuLK0R+VTr8uVhQmekv4PyfNvxgsg5OlDzoItNsiVt0
zuTWlL/Xa3MUjjJhmL5G7k3kC13CezuhHOPbFmBKtLPb9KlKFh+TkH9lO0pbWBPUJ7r8xruVOgVd
A1asStEvhffOOZ9ZmQ/yGO5Ee467WCiJou5+EO/m/W1MqPIJrPD/rlN0mubn19O0q+DbR/KYElUu
a1il7UkWQ4f3I1RayHB+mMabmVtpXv3QIaGHPjDpTPSEQiDXy2vMim77uv2NfYz2eGWsPL+ft/PE
BC31Q7fdNnJ66ci0M1Zoq1t+D4rXSdfHqTU0Ea96GYMkhY/sqN+tAYvvXkzL214MOk7f9UJbjSkW
zayNrEnIjmxE6ZAA1na0rbeBMaSauBxvEG3DpQUiQxEhMyViyrg3yUiIutd9C3ixYX1AMuikbEKS
DBLpFcBYMnOEdrTj9zkwg/ipuUgBcj6siB3YcfdBB9g4a3DOEy5HloMSo/3fkyOhJ6vX8AleV8oL
TWHS4bXsDYZfs+BiULY7DoCDIzs2pIhEmdVx6DWHBd9DSploG3k1A2hFcP51cR8YwsFPv78JFadX
bOpHh/rOEvAHJm36OTsu6Nl58l/5XankH+MAKMQHf7mCJ0rnI+Zt4PFbAcP9S4lZUW11BRuoXseI
0iJsrFUyNd8tpHkgOL4VUd/8nzVjQaWeAp62GIdtc0ioXsjjLe2nf3l+MhUxXXVldLkj6JezA+aj
Pxre8I4nAje2fiS2ql6z11AtADdoqFJPkj76bpITpIRHGQ+7vJZ7mwLV+AsqvMBp+17dGNvL8zFF
eMJoZG9AfXFx2pS8ccShiwzUfW2ws/l/TJYADVYt56LVvkk9Xw02k8df3tSSmo0XrGv602owNvgw
DfREGutd4Hgci2FAIABwtmCBFSHp3sQVZmvTAnoK5reDo87HK6AEM4ckIbk3deZW8qm79tBVC5vt
tlvC+f1n/rzCDL/f7tHPTE57peu+U/uVTbSdM8KosToDjRxF26c/qukODReqLnnsLyEOh4jwOmHE
hPSWYiXI0S2GvHwjs81bGrTaSqAQw/SIvbzOm9HECOAQu6t0RedASQQW9s8IBu3IDJGJIrflkIsd
V0xVwkTnxYEzBQAjLQWGpzVLly0/pOYxq8KnOGczc05q3fyWy4wfYxDa8LZcH/t75ayk4eWYiESd
Vps5RYuWafXjIX/qJH8PPeSogHf88tTQAWF3+FOR1T/l5PDsVff8AcvOSiaKbDFgw8B5/mCc5WAl
996J0KjNvfKvYuc2G1uhtutIgvMs+2VWOckD8qRJ3+qjPMjiK+mzn1aGME75KxVIViaT3qGKBTDp
FsA34XREutUkwZ5k4+n5fJAMJg72sW1Wi/lJPlTLYmX15pFsw8J/MOxaaW2G9dnrSItzOVyteNaq
6jNvQhlSh5YRWhgHhKeNrI5YFgPCyW+SDHAisMhn8WZJ9oO0w2L1/ojJ0hhR7B0iOJfNxaclylmf
nCQhgnvfKoM5GoBNYqfJET0uxXNFqlgCEXTBebE2f+vvysSP5G5vKHDJaeKSApy5/7BufNYP3vKT
iWATp1ltVmqYyEKUEsfdGC+Ijih8SvRHDRqGvvN/v/W84dtnlIk9tREQiKcD/bpMIvF8RhCxvdDg
1N2m4D9PgjhmmwrB23O4M8e/pIvP7465XLOjlP4jdBsnZsh/SJIj+Yot2K0wTj1mxKWpEdYGmF10
UBeqbc8jLMOZEsWgTLlP37iLM3fyc7pQMUfOcE6xqFsNlvAOlbjb7n+jt+zk7JHialkdYlSJkp4s
43IKREnBhzZQ+BKj6cXpUl5vSfdSweOkuvXMB0pXGB5wNv+hEttssoLp7GaMxMVBYgNtNalvU6wm
9CWF9QS3Db2NdVTTlWm8YyDpz0zaQCp8RHD8GmySx0+/5I1OKw3c7lKckjmF60V61xpiU/iLuu3O
UeqGnrwyXOveUu93TK7Whj9Froi/zg0wXWG7OPbGZXQ26ERLJ5b81/7372iArcSWUSXMBicCG0Vy
zvcsq/CSpgaz+VsgZ1F2teqi5Y7dqjwdUCKRhHRp1q250XjxT3zT7h17ZJixtUZq5wXHAutbnqR1
hnVAoKRgBMixQvL1Y0OdQtA5JYkVdAOW9HUpp/5GDz4JbtHHDO7zxr0OCytK4kuxgvZHl8IM7lWj
Kw+4bne/oPg2+qFPMKNjprP2a62jqORMCH+OgOe/ozGHDEoPORcYUJuY2mklH90GzSyNAq/l/WUm
ftH9KdIBpbfxEbNNcSGkoq//FbSfOjf9oM3B16Hgu1JO7L5bEs6qCJ9xtA9X5utaKdtjKK6kQeQK
jQG7mxIZJJnx/uX/qFB0adjreXepZQRALzTiIWMVi7UBjxbQRz7iOWYC1koatUivnLUhLD6wSpr8
02tnuIqjIPMf9aqpb8L0Anvrw77bvL4TSdNKuNAwc29gDZDweK5frsMav7nzvmkPGTlACGlF+1j2
r8yVBQpIEofSyeQJuQCqrkCjf9vMfZLUa141suV9nDz5gEy6q4Zu5ruIlJE20jCECZf93Oehvmuv
VeaJNK0La6L5ODgKJ76J/oyNalOYzn8ZoNdUWSZ8kC6Y8ObTbBBotAzbSt1hv+G4dUtkGLv2J1C7
MxrlkCjsrR+Gw4DXNmUWwiilq4zXvTY1510RTZVLW/J1n4NDnmMnDsTSEFPvBrxDCoarSeqRfuQd
Au4xNsljUO62A7R/Li4tgdVrbR4QBU5V6vnzFMFDJKdEkUtf1QuOf5yrsND4t6OQJvbYG0eIXtof
u3F0ATjzRq3jGjKaz8BciX4/6lq1dTrRq7Q1mTQsjH4MZPK7zL20OFXe2irr2oggn1qVztbJfIbz
Mdrury/hZsDvhcYoTk9Gnahql384lcK+UQ6Ij1NsqXw+T24JkwX4uwbES8pGDgfR+VWfb3+tVcmv
SWDZr8RNVczsfws7YvJScXwbA5cLqjINLS13G1LgE+tLviJV8n8aoLuckVkSF664Z5ezXtzC8t2S
PUGeMBOqBsfoLfcBX5aWUTFnCvdbmXroSrJzNm8IP84k+HD2RvkoU7JKUTbDQKbNBhQBRYG+hEJ7
tWbai47w5jEdBoVJSIg6xcIY0cxzjH+BzM9c0eJP6CqI8tbuxWVatRawKtNeCrq2VA0UCFQ3crrN
VfjpsTjfanFG+q5IeSVSkVWS6r8SrtWFFfs9vCFKhvag7tvZqLI90QZFHa3MyxuL7xDbY4H8RHud
ibwDKPC2wg/mGyKkQo1XOpuivUZMyxcOGleIm+pMtU+mqSJnORhExoRS/CIXJjZIiLfIofzAUFnl
LCqUIZSmjXtXxYgbW47UyJJH+q5ERHEwRocYLkPeAjORPVwSu5Yt18DVURA17MW2GkdHmTOO2b08
Eh/LW0QWgCjAr3nvFE/BytW9AlSQFV4AH+T5NOeRGtSjIfmzgUCDso8DoiT10teBnHDzTCa5prZ1
SPXSvAglF1X791qfAsQTYG8y3xoX9ior4V+VI2QdqIWRal+dUs8z8asWJQE53jOfGjLDV0wzPX5m
0D2itHuK6aLgwyeg+fQDnawyZ0IHvi1lMvLwLc8GmHGbeODIqY1j9fm9r9tDY5SojnQtyeuk82NJ
dLIpHog+Qiopjo92VsdtYywSuMtPLMCDvBajFG97VrwWVoH+j8CmWaVw/zmoaR5FV4eLSnJ4ROA0
rcISfNi+1Xma69xN1Yu933/FnA9jdpSix3oaIe1uI5Iw8E+6+RwHuJsltCjw3YzUg9/TyFd7M5Fn
0b6h+p9f0eAG2BZVKIFrfXy9HRSjIjB6/G5gY7xnoXIVJD4YrSPlbgcy6AM1fon+b35GuLz1YCQc
83OE1XEqHblUIXDqkDZu4EugF+6kDmF4HQcnuHa4ug5R8SBfG6A4mTnPZHu4JBxcmxJF8FLUbG55
tu3DtzKCbMoKJPwqGH53P3h8JqPX/Qqq8uZ5lxGeyX3D6OtFpCSkmlJI1VaPK3srI4XwcOjnEjHG
9g2VssRXVTPi+x3DhlDzMjiXg8Mk8/e+eWF4VE6eqD4ZUemcSpsdW+M1AlZ1yrzn+J0Cs9THIDCZ
pXPh51aw9OMF1usrM+eyChw/u4PT7urA1oEb7ktAWNN2Pc+cUpir9UNNZbhYp3P8hXhqntRlGxp3
Yzmm08bqiDj9p51lcor00pzpaQiph2l5F9lNbqrktSahYrKXkOangBoyFFs2PeBQcTn8B1itxUxm
+cG5wd1p754/KtblxaN9ynQf45WuEo/vC2D48hZNsBa4uPsIKyrHoKfePj74opH6Ngev3JN64SK/
JsfzbR3YlW0ozvVkF98sq/Ett8+WQhSLV7j3kpeQQysKCkjESeWX85uiAcuPaREZu3FEf5ZhjF2n
b28Rx9mXSl89mx0po5iN+atFYWnvF4yuAtfwh7A54Jj3Rkb2IVsm/h1fuc5HBOi49V7nTWxzJPZ0
ZaIcvCLbGSxg6/pbzjUzcYNd7Hl5hm1Qyrj9iktJSMyGg4B53dK7T2k6aSedVCZMAGb6j6bcSdk/
XBC44PQQNWiC1lKTAEs7sXFUt64UIVBgaBR0uPrYA/Zu8aebWEC1xLcQz/Wln34phECpinIqhUgv
MSgiegzN4dzwSj1AI0YaTpxU4YPLxiWROwFAjrUjxT1IOKOelqvVCUV4RC9tcqmVdJkJtLjK2k2V
xrW9eR/153bSDsPzBvwHOMVYVKc44zg4oVkD5eeoAGSncFUILY3s7jL3aDZMtI/cOg4Op/8mRDF8
NOcvjar+5Ko6tuUc4h8xjxN/s4/qPAN8wCgwoc0aOVY4fglJKzVWVGjcec9Rgpo6BH1Mc/6i1bF0
K6oyVBXJzTcr3bAi/pKYOBcFJvfQbhjhbU2GGOCkEMR+eTAwIcUEs9tJz5Q7TJ6lTkBnmH5g0NCY
aSoJs/HO1tSEqYBFxlIj/vVQnK5mcfT8LQCyKEGDH5+SQoTXjEtFTjwI4p1LuvrAqx+jGYZfkwDa
xDn35ZA7bXhulxFdmemogvEQx3pwLuPpu+YytDS9N/9wPo9Bz2sL+f31hwrylsqDmDLP330I4wq/
onMFebPn9Q1Af1FT81PY0AE2eT1lcjdyw9sxuK9qDWjYCi4SX+dbAcAOb+og8F6UWOqDZlo5SUTQ
9IPsG1O+sEcDok/XZZFsoTNu6nzLNtRlNmWZCzzP9pbCsOR38PzDqr/5QDV1JSiHwn4LXXT2dXdn
VziGOUKMhrNG6qms6hqQC7gYFyaSZz0tZbArv0a1EnJ4NXQ3aF12FDJ/o2ZG2gZNwhtJxcO5jlkf
wfVm6wZflxnTVvHcilhN2GeAdZj6sB+hqZz4svd6OB2fi6kMlSlkkoZaB6S8Kf9cOr+C9JxfjH47
RjQ/3tW7pkhc1lhU259b7lSnW1O8CrKo6JWK/Vx65cicUrysHYhbpy0pT5Nmm+1/ZKRAkIIvlAgp
aWLh1hfw/SyVgh+XQYBevBqhen7jtqsoyOmlge7x6wjoJjBMYyMnAnxihbarWgSezoNmrSKZwuEB
+yfol/XoqQ1vNRBsl8SOdmMHhIYZL27iDqjrcVWkI4rCKZlx9nUtfreoRxn4twPXbLJZsqmy/OaK
Q2Xy7Z8iMKgPJect3zo8xOJue0IMcKZP7m3D2/7JqHDXLKZ3T678SVf+3XqIxbzdw0zqkPjOi2am
jk1Olh09rhihpvfZaXaZFcjE/Bk8r7AsL2nWKf80PTfZTzIXAEcslt6rTDPRgIHjioLkJQPTPM5u
lN8fUJ5UoM3laOFYtIAKtHKFctcX/QRhcWu15y0AY0pePghXq4jTjPkzAXslERZr/nEYY+cgV8bd
ICKhH9LdhiU3cYmKog4pzCdv8KQHkCg3PC6xT1yPEhOA23BMCoRFNu5YQK5Xuy062jABz/n+/NEm
oZTQUiegEpktXEDv8XD9LTQcXh6UWi3ncYm1vkIey6zif3lYrgPpw5BmYnaeRdgrP4gUOfDpg4mc
mrTQ1s69okRyEGf98KGDaWCGnoaQMFjRC8no0B9nEljtJ9pb9GUMP4pNPa5Wblo0wwu/NNZ1t7Dp
iIGpSJC5JyqgM75VqQRaXptBSCDjqdvOhwdLRnYhl2t0ZeV2Muq4D9HSb/COdkn5SkDWTa5XTs4c
CH20QO1ewenHCpKef7Ztd+mMLo3uOWXx9T+ePOvRDOwP4+mrP7LntLrin7ZyBQMknr72PSAlQB5a
4MoWgTKMdeEthazAgx/zLIm6OIXof+voFlAjGs/bfBpAqUGBWGspfQ/65SO0crY+O8Gj7H2Hnn+N
8+DclVqnFXvM25EWTknWu6ru/NjGykp1QXAZTJbzwKVUmvbaLeo/gWk+FYEbKI5PWU/aKGrlU0rl
RU2QzPCFkXH/itlYIjPmMibo85j542shTFZCEtSuFbLb+ICUio6BvdesW39U5nKgJZUXlYFdM5xU
0wDNBEsc8G8CiYgNxsE1JfQkZEjezibK46YqabXqKfshafLyfksC0hUxTnDiF0Jk+SACabdJ5E/k
gp+AKA8coq8V1oad2UROFnkZY+S4SDPltkSGPQFtV2WqrlP5rgMZGdUWVfce/NdGB3fgVMxiEGWk
z4iMj8agsZwik+9Z9w251i4WreuwhsqXB2Wc2ft0Rn3i60ED6DmkeGyUC2RW9qifaIgxSbSrEdLF
NU8veh3rkIaIXY6jBzB3F8almBLsMvOoGB9Dgame4uSA6JM2Y0GjurHQtNVfguqb7XundDXSgJpu
jN45oojHDLqUQEgWQiDfTSnSviQ8PLW49OklqYKwXoP+hoc6rGKhd0+jOAYDZwUN7+EODpsbiEu7
G851sI2CqRBnBtSnyv/OI+5/cTrWqNPbhex0tZ2FqTLzaVvGd5rCUodeHlNPScfpEFP4ar9VucYO
oxa0ahqcZgz0p91fwu9toiettno/eH74uFA93jOGcXglzhlV2A1fhcZE4XDag/V8QP2s4d0hea/8
2XzPY2G41QzvevHDWMR+quPhK54gQwWGd8xeSxd9PJPAT1tjDAYYQyZICjaEQ06DcLgJI8rfm5RK
T33hsccAhhA/8COfXEAT7/1UjPjBHan/VthQfPt4gT+UbR+LlD1ad35dgONrQS7yrYK/1uRGnrFT
gMhjIOGYpSBWxOYzZSP/Iw5R4HS7Lc8MWLjdUcYrLR8QtRP+nU/aTYVsZADDdvqZ8ncxS7Mmb0r5
Dn2FHk6R2pIERCBLh+0/T2vIecdL5CNb8pdshjrgFSdgJF4M1JMgzH33EZwNlQ2mkkHBt4xLV9YW
zSxsqhv/a15JxK6PyUotaj6t2gtx3n8pI6m+eYDTqIMTfnZ/q8jqczJS6Uw3TE3PzWHWcREJL6hW
wPeTsi/BNOcCTnH47RWh+HDnAxseNak2KPm4AVbTCYSM7qSBkAp5/zBlayHcGB+nG6MLiqQtKiw2
JmTEMYTzKxGZISOCPfl5HSxOHH5C14CnE2atmNMqc5EBBwOAVtKXLwQufVWCo7CME5FmmXC2yTYc
qBDNaFZLVAUsLB9mk+aqw6c9YdCPIpUT2SG1z6O4QEgI/B63d6gA592urufMAbcO5e/tvFD/qaIl
Tuc8fJI0fcbqzJxZIx/yUGTyS9+UlBXGBjY8D3v9tYWSW12kQH7tQO3jCvj2P2DqFX2bMpE5TrZS
1zX9qtcM5NVzXfR5FLB5kXLHbFYHrKXhXg3ShdPQcHpACPPfGcW0SN1Nw+89HoDseiWS3CA+LGYU
UsnHsZcsV1RkPaH3LlvuRs6f3CVTmnsN0/i2UYt+j/oznvLW9GHHZeDsJj8lr24z07zo7hqe+i2W
Vf/Fv5kr3kno1+iZlkiWGqr+ZJJqqil+5VVNsScJaFpvgiYex6LSHx1V2idXBdDMdui7RlJW5Z5u
caIoNZOX+v0BHg2F7HUKyT5G8byZEadaZ0DptoAl7qWCxB71NcCZwtZ6+njmCydq7BvfIfg6g8l2
vRm3Vjk1qEy7K49/DU9rTttsKa6W/8MObgQjACxRpVznoSZrQqRjQxUrPLrbruhv2Q9c1bJMP1Tb
nwds6/PbS0Kif2pLw2dA7O3rWzUdGggS88SaHh/3VjbDv0vvkJ/NcLsR4wFyyoUEo7qJtPCouFej
n21BJRYA3M0nEKWi1ltI+JpzY749bY8iP/t2O44kWzFPiLoDw/lpgfyUZVW8y2vhf+boTqGgOaOf
VF+Lb/EOY8YEEtF3Qe6Q6cwNWYXS308/HsonDVxcL7LXdfQDJRsKvE3JFDWxEqFkKO5iBmeXP5O9
2VZAZPfyOrwrNW3x3OQn1EXzRWW9u1rt7YB90XSGfJH5M83pP/bYrXYdt+vXoSJ6ocAnzAMrpfFe
N2eWmZj4UPci8O6EByi/fx2y4JCNjUToCCttGyqi4MulYnXTWm8JMe7IHt6BzkvcIjJvtPKKdZev
ifNL7CFEtBczRnI/8Kid4CDcBiD88NrLydJEfqY4fwqresnD2/U6gSGy1/kwBze8LJylQy9lou+h
2c3C6TK8PYDSACyHcBU0RSSG/5M0CZbtPzNaY4uO8k5s7VjkPXZdL6bKSxSyH3I9MvsyItWmw97A
dDUZysywZ6ywtUIfbkvr+m499NC6wyqvZTRA5+EdwDnYExRDWGldxSHPpN/gN333uLxEbd7rLPnM
mL0hzo1OoowWeKkkFrCFJSDqho7vN9YHi+JwKjv5x1mKzozTPl0jyL3DMrAZPgs0KYPskNi33QMU
hSgA4rC81tUNWSOrwNigPMLE+Ekl48x8pwMan8EuG6Gillr5ebIK9e1GhbnFp/yEbjw/lraOGNF7
WQkEJaVGtKZyFISjRLGQzhHRDn4JcsdeZri4CRGBTRqIoMsgJHfd0REUBJc8mjfdAVjVwKkIo5Fy
GvnlqPSeewMlFGZ94eNDGSN34s4s0B9LYjEVZ2tWu1F+e8W7bCenMtm/3pGVYcdrp/s4fu3viiKe
A1nujArjN4La9UOe0Sx6859eKSTdCLSjzpu/tF5S0Nsyz3889u6xVO7+D9ARUFhUphveiBJNVS9N
0nrDExBlCkVRBT9ghZcJAjCE6wRSdTu0yoAr3gqtcZGjGDh4Q8tiHc97+CV15kJCjVM3MYF5STLb
6RKebNmcPE3lagTeXfIgwxecuYX2TwnKaNNmNEZJAiPp0UxkOAFU25wYLpKVB6UcqHyduc4BsI6A
8x6w+XlvvdnfLfJonnkGsPHqCVNJyqA619CyqSZV4YaPrvHTbr8PNT+6hNdunXTFANHnNQSejtVa
bdkf9mOZhmlBon2+Fe0XvmBcscV3fRRmFto9Rl6aVGSGjJKr4IENQFAqHJk+tqMs0vZf0trQOyuI
ImHyhV11GyYsTh8a3Hb93qwhTD8wztYbbOQBQSNMMllsQMJcmsPby3Sxl7bHnnoLh8lV+PpUYrm1
CMdmauH0u9fX8zBo8n1oyMhkJ6u9QdNkQkRRxSXzINVo+OxNakeCFdHWK55On8XcoqiikcMfM5F+
St+qza1u8nsli1YEuv/0XNBUhkNwG+Vr4HQhuX7Ycz8DvesuTocpZt/wB9jVDNTV4hcc2yrYi7im
/Ri4240tOsZ7IrP3H6uqclqoqfL+rSzEbifR9km6jZ1vPoIZkuoSy7+kXTZM2Z+4ql5W7NkJz86S
IcWTfPv2EGJYYMRCV4KlK/Klo/XzNl7L7R1JimBx8ZZ/OUyHmX76loXtatcLn+ABZVFty/eZeldq
dlQa+RtP12ViAns/4kL0SiBr3M38Sxl+M/RA94MHLpZ8zcEVzSgj7Ep8y0hB+Qt2Ea5mVQPvlc3A
b12gFBe6TRlH9bG1IWURh09ms4bjjUitSBms26D15VsWPowLiEIlHNScV9uVyVkSj47a7vaccmF6
y+4LEv9MBMkJOpK+3QmMeUekWrHkwH+T+u9hw8QlddumV3nTvIBQrjLM2aJsGScbqNGgOeyup2qt
kXV0B9Q23ZOLxrdSOnByYJtzG3Mm7HkP5kLVDdfVn18ATWVXCqxYDFQDYBeZcvcNcytcHEi8KAgP
Xsd1YAkUsZHu9HQdlrL9Pxv9o8La/wVhOxvwg088IRb4f7lJQyFAJ8Xxnkp5pNU6ERLQHeR1x/ZG
jiJoLt1oIg4dWyUivDW5E8e3v/f9lqo0KMfMTwJg1rN5MAzvNvxpSHlbVSVd7ZSj9L/Ca/6yCYFf
pRrULQO/irqp/Jkn7+iEjnfpT8nZKteUrJvK3xmNW04cQzsnsj2v7sGzw7nOCqh0vIbxeEaHQUmk
rLEVEO2hDadyHOJATWKFnmUte6MM88eiIrEaWdBu4j8YD2Z8BW30G8/imEcnMtR23OM2SsTNGKc+
o3CAMZvaCCecDDLfjiAe0zsxb7htx6HRFt10EIW55h2IKpo/dCI94AJZax4ebiuvuPi1hrTO4zDo
vz5qpuQdA4UpVdyWpm+ON9q+vygFdAT5cuutaUzvmH85LWmg+Cm85sMkwBs//ZGfH1ihLu13CI4P
jlaot2dS2fuyuGXLU+93fD8kyuDy56cAPwyhG9UE1nBzw3KBzdmn7lj1/SRPE+ByheU/I0r0Su+p
/bxfILFdg7ydfVSsEigyuIdXEISjocJl6ihe/eQVSLPHWxZAn0ez9ml+oSDQChL5L7FEIpUJK1sl
mqb86k1hpUkGVhXuhdd3WFKX1ig4ioyYyDsJCvo6wcinZIBy/FZPL8lGTDXQ+AGKUOK0X4yrfynS
+zQjXx6PVw2KFkcVmbwDmfPP+yP6VkWClSZWLTP23TwWK+qdrnWq5OA0LsxpuPGhwrvdMQ122pAT
IPnt7i+BK0Zj7vrlTcObco4fujYCsecuXygKT7q6rZwjLa66jYef3odt7gSAQ6eWO6B0Xdkfq/IB
LLw2Zw1C94v+anPQnLs+XddTfymjsUnr4tZlTaYD448aYgHCgcIAPQEnZ+w2guP6RuemZL149Eoy
yCYPe+vkQSkqKbqvYH6c/49ehbGrgl3bzAeF5T1SHQfXBzjdGIbHmGrLOlWkIu9GjYJ34SzUIjrK
fJCStRDp1jj+poGRtV5NxFdEwBl0FYa+DUH/2z+qhWkl/dUrSS+Eg/fAtyGS5ERkyYuKMHeV0yKL
/nhE0BH/DcN7gR+hbpiJ3Jc0AXBPWFZJXkCuJWeRc2h6W6xDCMetNJtDOXVI2xiyCNxiGETbKj7V
/mwf1U3tDx8EPT57B7PaPR71x8mhPmWLmyu1Dc5eGiTrSSICzUkvi2ZuJVa0w4z3y6AXosIIm5Mw
DKUUoEwQPrh4oT0pPvWT3n18cYpBdrvp7y7GkASXTJpIijCauAExJvFT0Ggg0ejN8YggnGAgNhGh
pfNKArreQZ95xx1uXan7AZBWRJnIvz/xA7xe4fzRkGeIDdnxKTDP8QzaLQGFvxtGHgt0NJQuqCFw
/nuejTsta1CyStje3+L1RtcXDXtqTggTS+nLlCCo0KAbIMbVQuIfA96lMl8X+53eg+owhFU6GRXr
oT8+RaOH1RLlaUHwlNPkQwCHpfb72h8BRZVrcg8tu1GeTbateziRWCC9Mti+WK+x3RtCZPwks0RN
rvMZ2SeXc5x9XNaZQpcJPN8jwfQOK/2eB+MPwmA3TG3jTDsH4H/Kd9KciMhGfACrDVIjaCoMU5R8
j7tDpkopLeF7JlNraQHcfHFLrrccpLduRl9RL94yRe4vb/q5kfEprgbF5u+eTOEBk/ngW5bzAviM
dR6iUXBNS+bYDoxid3o0Rmm3wqHaNbOt0RNgnLM18Ru5Xk1Yc1tMCxS+OVbd/N46tiuDZmsRF0Pi
mMgGB6xyAXzBqkJ8wv7wbRPB4vHMkuiFD2gYFQHMEzmbaSBlEXBs7Imfv7Oq4Khxuwqu5txmke3b
G5LRFxDBtHlLaLm6Bfu2UmQ6OIWL4siWdDVKl1pJHkpfCQiTVy7Ck0z2nRlrNR/S7tkgo+WpFNe/
KXLhEm0rYGWR3CyuBIU9WWqDVuhs1bA8k19rxSaw4ye5HSQPcYuP7lfk/KqHFfF7HTVpY7qYxtk4
HPbE/5DuQTpj8Fm8SqIS4uRA7x5NTQhZ9/a2QciDnuHYBbrAwU8oJllnBpEmBFxlC9KOeSsOWGkm
6VNrJQE6tZwcWOOk3tQhM6Z/jRmofsjXOZuSIcjhMuKeyEMzdJbZ1tkf6tcnHh8LmJS5tT7ZXQDb
jU/EexSvaZMTJjaz8xVj8V9V/IVAULmYIdUb7e9RKwKcsYIEwn0y0Y5mTIEnY1jJ+7k3v4M+qgte
BFLSkcTatyS1H1Gdt5ggFKSdXwIQA/owWkC7dXf954bUvl0JOXUeSu/mYSIQ3Oz7oE+cm3dLmPwu
F51hPrI1SuN8xvifbybsG4MEUckXVJKcf2rvwUqitgSo59tjamSIqTfUOLXTz3HPEaG5fWOunyOw
YgdcniHh3IDV2apxxCzN0CBl/SuoKBk/lOy8T5c40X4HL2+pOvrVwV/KIQzDA5JaII7I4GOORZKN
WVHPfiL4e7+WzZpJBQHBqjPeDmnUpg9BIz6su9S0clFpI5IEaXpTTo5ywb2nK0T7oXy0VAuarn+N
NTwHdYWxFPrChmP8EDwXzjSq2duURCuGo0lHz6FknqoZltwdR8fGGdO5SKELSa0p/KY3Rt3bi2BR
8ip3Pa/2yBYoW/Q6lTWnsYrgW1LMFAjv4QxFyKtbHo1O+R8yZREaNFZF02z/k+VGRXwcZcs+PPxR
ykY8awlbc8zw4KNB7wxlK3TF7IeI79RDsbxmBK8Qfc4Mrnip/ZW893YvOAY5qY+LnLpkRAQNpgj8
DAI0wuKBdgPc1pmfPAZTd2nP692eadkxfwec/NfDb1m/6XbN0UAMxX1BDHxSKfRCMg7gsKxG/qPp
OD4//4wtIs2c6ULVhL9qwsQjnr7W1avwmVo1Paovf0Cbufl/Nu3C4ykSlJHYPyj+xcmRMTEHIV1y
GV5VL/wgQo5LTPWWlvnBPF+oOYSIe/YXGoykgAS7/hicKLPXFhYe/Pme9K6hQ4IzAJZBbEhe3hLA
vWGSZztHu/yus9ncD6pJODZij2pEb8Ea1RGzuhV/UTwIa1XrbepHiHSWIi/xlavI7q/EW2QB2C8a
sh0cDwdshOd7J/b9bKoWUCxXhH3XFdQ6MGRIrFGQ+wEUeM36ksZXRUYHlr9iNr1EJKgABe/YJWX7
A9UL/6JJmanXKI84RakmmX3vxoTaLRsviyV70OKcUCtmnbIBrxoPyC1ZX1rTuS+eD0tUrWEgdqAg
dhpOBUnI6WEm5CDWcQLq6YCk6f6TOhuo9u6p4IPhTY4/be2IdmektssnEH2mpOmCsPh4p6b/9A6R
MlPD3R9lvez+ZjXnnC1Na5SceVQPxAzOKfaxDEa/+CoPM6NeerNJGbP1odLNIz46hchfGQJvJLeC
fZyLW6+N4MRMpzjcDUWkkrRHWa6hrM3FPoEQ/sbS/W6A2di3v30xYsduhcmVw9Z67E7eSPoMwmbw
tNNPyaoHwLSinlEzodQCmqNdsyolaTYvd/8YbL/nYzw/vct85FaGHIZPXLaPPr36uMDzQgBtI12+
zBg/B9JJKejFpg/9kHolgiXed9oP3VI5tgS2iXnqubtlrsmdX/dL4mNDUcTRTsGxFIHOHjpU53Wx
eLMBUH2+HIjoYd2QxiDajPWLLyMFHqcPuCpxk5zzksaVrnHiX0FTuJdjvgcKhcIA6vpApGjEa+ei
E1jviZy/2HrPSxddShmEsLZygCugfayLKXOrj0adcDe58gNF+52sWf8k1VU2EUoifo/1D5yXqcoc
ZkXQLwTZmIsijU52JcCq3dITejjr0ZYqV+3uJnNcUf4g3n2fpgTnfGX/JDWh0dNLj5PLwSdFsHPO
1z5Z7dr1bYVe6QItoCx/CqcqElseIfSZJ9A0UX8SW8Rox49TqpYtnHJU7cvEqNvxt7bKOPS4urH/
E4H9h171t56mtC9ArXLd69gNMXD81twePWnzKk67lXVpVQfNcYRnfsHrMqQtYVZAdrwWT/K/txgX
13pSC/Z49nPKFLVVBWltbHLZyIxSFOyqZiKOXfjGFPlI5oqj5hOb89esKJ/V8bw2bdvRWQcZ7/sV
0idBhNz80wh7JUa77y9/lBIQoivZc3tTL9oxKTDKIZ/+BO+1GMQPKT9MZLrYUPB/4xXCQKeH71Ow
hFHVMQ+jjVwri5dPjmrUeQ+C+k9b25FQ9n8MKcrFygM2rYLq13i8W6lhmXo7+TPcjYt/wjysKAJc
VBfSX4KCuh4+PweVvbptK4D7UyLLDgYjFGPYernmWPu3slzfE/MGxkeLRcfY3QxzpLTgMSXfbKm0
KI4pW44penr/Y8OVg7T1Xjp4jTqwQYNWwkeWqG7/HAsHNJ3c6Uku6k6I72O5H3HNvllkYpdjkndc
309ChQ9mYHWGDu7Fg4J5ucVgS7SUQjXKkN3pfYIPWzdkGUhdSyDvzlTAr9aoJakBlaLBZb/35m29
AWJv5IBMtP7UEwnI2JBcC7QrRFKfFLeyqjsfUxUpxv0ArtCHxiiNWMCchdWxSdqnXR6gvxCi48qo
4Ug1i+q6YgNBIShSQ2Ewi2R565JTD/mJ8+drBhUb+uMsWTZtHRFj7ACqtXWeOoXfn6T1dNKBS6OX
jDrx4krRZLKYmbXIajJ4pBd3I45alm3gJtBiYAntqbi7fTWvZxHNRRlBwLbSSFPmORfs2oKeghVO
9DnFA/rEF5UcpEhMivdyKX8+JeIxscLePS0c1byc3yJ7dcvdlH8od7dag9AlwzoATYVa+7vMA0QJ
0k7/SyiDwnt2yYg29HfEolqsIx2Z/GxeM2du0ZDSJh/yOKkEMEbJ3ha/t51KXAmwmTxgyrTQY0CT
DgKwNiJrhCcDpUH1ZSdL/WlJsetsqJX7CialzSkYD9xZvFL6u05pmS+IIHkBHb7OeKIRpNYH8S5+
9DN40n6qsbXtxH8Knzarx4p9+okqQcyg3N66wQEv43YQ8NzdOoA1fzDgAEbszfrDgLx8WpCtxDHM
C+NraK8QuWzwYoTfU9FzLHyXXM1mw5preWrrvYFHyEXKdos5BCDsS2AkBMV7H0fBvP3/ROcgk5kY
vyXmTmCU+QgtZ9tfHZUfEdgemfcrD2/Qn2xVKu7bMyCeiYGdTZwvCcL9pFkd20bI0zmBIk9LVGaY
VbMmubbi1vz8Auh+pL0NgHF6qgFnMwfySlbS9577TUIiFEJOEQzljw7MF9YfU5QwoKSnnWt8o1rC
/7Mhvi56aw3PnYjCMTvvGoRnL2Ut5GJjst/7tdev/2dV293TGVAespsII7sNFpQKpkcm9jdxZpW6
9yvZB/61cybAvHcFbQq4sG9hmo9XKftcwp2lhPYssVpVaailbHdsV4mMiFTPAbQ+zD723qVZQ5cE
Biq/X0m/RHByCM3wp12BY6W7UgG26Gqjp+L7G70QiYdLzsmxcfSjES08wJ1gLUnL1JCJh/2iP5tJ
x+e/NbjHX9LDhXl+uDizhCKRE+hHW/WwYr4FIKWUSjwXre6SV5lqfFf+6Iq0THMt4TGdh0TYeVCp
SxQOsb5Vak7fm2UxuLMbcf1/agW2l5snvDKQ1xFsgl/no0euWCoSkH9ATEYSmuDoq2Xge3MIAMC5
AfqbzN3cK1V5YNQt+vg6nm5t3FQuTGP1Ho+ETqoD6voTDwGruQ5iSEuv82usHjB3Tsdt0MsJfDzq
mbL9keFlEk4++2s+zDabOf2jHC2tH1v6q5ETXqQThHXBJ3jpf+kfCoxsMqtRpsbda391WKNwBn1C
Tx9xXXy29wG2IEsHf9BlN3j01oeUrnr+7zPt8pRhRrNjLWuWXXdOsyut1eY+nguWzVPmG9IjReuB
xj+AVBD/wDqN+GJk56Tpl+Gyj1PI+2xmsKFk+5pJnQ21WQZIpZubMHYqX+ULrVF17Bp0FQgcLjCh
kmWhyXIaFGsJwi4Zi112DqyZK71gB3Da3nQzjOvPUvzNvlHSoE8igfv0n9eBPNHESecy8Cc8wGrM
hpenlzN6+6rQj6IV2hJYolwq4r67O4cwT4OtyoGmH2C5bZXlG/3nE7g1axqSWCNwc+WbLT3B8wuF
pBfCku8jTU+bikVsItUoIdiTinzwt/7pchn1aOIwNUIh2jAtc/MvZfzArlowc5j36FhMcMeJvoUT
I85syy6uzBxP6d9byOMykGIba5uxLuIJgblPN+qzpn11r2x3YkIr6Nr7zjOmuOdAzlpMM5lHzx4w
+K/Yy7QtuaWzpbzSotwRbZD43KdURxxA6iYZizNaN7aBUbrrt2gZuMPDfGg03CbQCz3FrC13aNGA
cbXdJuWr056Y4YK8YZPozG+goLImqy1yKQS7W71tc0Z8PjOmdmxk7g7LLknCfiI1RSsUYXsFrU7s
vKgVNtv+YFReHTWu0ojHVtgRIxvBZk+bZbai/gg4u7ymQc1Fd/3Skg5guKJ+u1OKWtWhMdN/BZIS
n5h0t6hkCpTaNM35LlOK8Qa6FWbVmiLPfAPUo+q19lVqwavYf1TitzPLL77F4Rs/JgEn4CueEk1o
xeJGfCAgxifJIg3z0fajypO9MC1jfAP9mMMhulX+/CROYlQFWtJV0thfTQJTugEsGYmIYOSa2GZK
9EqlqjDjlpCK6Gvyrg49dLhObfZwJ8QANJ4cIuWQlbQIYPSmjRu24BfCu9/nF5NNqJwWjPjXk8VK
KaOvuVOn/ijoonkT7OVSXrrtAcff5l2P8GYvCi80SvkCKWZwP29ykI8c1srU40iOZlfwoy8PvBpK
2ONZxeNG/pwHM8s+YmY5v9U9yM86vhEGQCtgbBg5njohKg0qhNC7jAcTihBUJSdVng+IHq62Ivhi
awSMsbbR63t/f7kXs4nZ+BX/0YnFsChaqH8+QnnEk9MEJVOtuLR2X09ZAK+FDYv5hQ1ugxcyy89A
rGuqWQiI0jG3V9tYe2fNIzt/TqiGPG1vlsrJbAAe2lF57v5FkcYPsL2bIiSewjmYKfRw3uKiAUOn
l8gnsKsA3Wg7BsMK6SZVG5bhJvEf2PsXalq5gGqdy4rkfPB/CTYAZvSYmcGfjamCkXi916jsHyAF
vJgzCn7QZesbhHa42yk6GORKHXljLHoNp36/MtflBAP2EbW1Dnplb0rSGjw1dnpazV6QbZRUGuZe
2jvNlTq/bHqRGVD41HB2bwfCE6pPP0UTKQzUmSdhDY/6GWI2JVz0hHQxKt+jMapvgnFHH0Dnowz0
4jz682avCfu7YTnccSg3Tb7MQcM1wxO+B9x1s/OwPWU31IksfLO+xy1DLddDIs2ZQRNilWuYw6rm
ZCid/Xqh3N3BhI98jEdK2Z4fsG40OPLFZvZ5Uet6QZzKy7k7xZa+6oNdPAZXq6M7tAz74SAZjLMm
h6DnGUzqG1uWl2EWTdwZ/M4xqkRKptiBObDaDULm7ogInN0ma5yZAPNzBl4JsEWIxuR5DaNPegkm
CfKfpkGAKK81elUVRcDTF1gegME3hmQtbr+9Ja0pTQrPo6YcgvZ1wX2nCjyP0z1OxpTHa++4F8EU
yq0ezCBRGc1BmIPW2+II9CTIPozTx/Q0yznrGDtfXGUoxxNgc7DJjAELfpvdlBmPIMgAaR3Sinzw
QBfhEfvDjoBlPP+25ro0X3s3UL1tduJPlI7ytD8YVXANdzENcYTt3sy7AdwFKuDVwU58gk04+Z3Z
gVmE5qOisDybDEzuVVZRhXmxjQ/JRIm/ElCpxMoeT+gKKMlvDtLTEhegTe02+dL6Jryy9w3M8JtI
0aZuraUWy6G4h8bLnUk3SCQBaaj9gNgxEqezubLGW9pFtuU5Nd8VFMlJkyQ4o6tc+pHsuxkcJ3xh
blvyvK11Iyy0UxxA/daBU2V0kYiwU/Af2y97KamC/AdDIzKexjpNFSQZ//s3HnLEd5Vtjy9ocCIE
R2383HhGkQxjPFs/e341PMYH3BjE6CTHQi/eXi2XiBv9Z5ZcoCfCztQ6hYJyRj6+/20hSi/6XuLh
S/7fA1ci+wMotWAEBXKy9TOdwwJMXqhQfCaKKVlNLDvbluW9COKz0/rSGd3uo8Hn0VlfQ5zf9pC9
+v0DcGqIvIfr0GyOen/l7rrTUAhtH2oQ9mUb0vF+/G/xd69LpXSClb9/aOQfqh9eeb0kKjhb5Yav
tWKM76Y/lYRI+580qI/IL4qli1Wzrj0JS0T+P2Q0+kiE5Hakh7tEUfiL2I79BUE8CmNKASyVUAUE
ODb23Z1uuljIhch0Jh7YY4SwQ4XEUT2uVJjXTJMrED9hfKej0axb8WxWBCYhlqGlwgRlOwf/8z0+
WGRDIhHiEG3eUtRwHGwQPcChqfqKjm0c27YKyG6yverRLqgLlRDCXhM7bxcTtmsNApmItNXvNNFl
L2ZnQp5HHjhjDYr8t8/eP5VH+BIKI3N3+lcI5K1eDBWJ5CzTVOPpryKdKV8i866C4L8C9T7VK/FI
it9hbUSS82Aa6DLqifrUS/ABsoDn6Nm58ICm8muCjzk1C4oCJOVVwuAm0ebfok7UxmZwEwAmNUX+
mqyEo/O3RvvVNuHQJa1eEPbL0CTNi8jKOop0gNoX7rgo5CIZE5PvbyuezaEg8WCkKVofogVRgx3b
khjl9vqe/DOYokibayJJVzbrrIr7XUPf13bdnplv/hA3DLr2wpb0shEe34GgzOW71wIOSJL2GYB+
MpjhUGCDjVppG3KFHEmHnuP+jZoQ60e9rbEOXN2tU20rySlTdlnaJ+lvlBONOjW25FRlAkf9jmfq
eXQkBMPOVj1ckG7j3SkoyBLbgFDg2QP7JvlxK1f4GNri0pntAzscQxazTX9ePDRVWM+3G6kjYwxx
Kz2G6aheKtzFi+w17g5cvFfkCkj5cGVtI5yyRpAd9psPWrdnLWLvgekQtEBqU0A0OsJJwMTNiIAj
VR3TlVuGs8gf8zCBo4v8E5VbrfJNEpzGngjmaBQkkfd1Q/rKZ2Z2TSXD3bjYAILVGAVjbKA7G8rV
ZHbO+0EbsVgGGLNTpJrGb4VcmTh4cxVTsvqmZUCjR1LLt+bh4dmQh2AgT4tmXMNyJLM/wwSm6z+J
HFGmlw1kjdgfVbeyTkVzAXIty50vzRi/UiwWsDbrgY5E3eSOx/dCw5Odeb7OhnP2FkaBM7w8B5HS
mBs69ZYr8jaoBqCUSsXd4b8g7trBpWIas0/Iw3oWhkjH/mUZQUn0FlExo1D6GXGq8w/g9EHFeaSC
nrSzbfDFKDuaYHqLYAMqRc8KPedYaQeXknp/6lzqdIjSlpZV703B4uRwX6l1wjGOmSRjmzrpXLQf
wo4xFxJFnB52FloY3g7gG2hAuPT3/CTb3DdP0jne4v9eKM1+CkecD1mgVzXVaz11FqKZGm+vLlxY
R4UHkHvBltS901PpKSljt3YW65AKQ6Qpbrppa1yR47+4aBNnWLYIhbT4/JXQx/AaQYaXBgUfaGab
7oT/syKNLY5++CsYD9OD79l6q5E5t3yCQ2uXh52vKZDtSfCbQRPSO8agOv3BDt+jkEpmt2tJof19
xbsj6LvqElp2BjJKBOfG6kFUwrjuf9Rz036W/f+lFYIZ8rj6urqMKaxd3tAIAxDv/4vyjvMk/eby
BAwk1RklaQaOlQ4io7cPny4vbv9z13N4Q90PbANV+KqymtJkmgRgPCXs7WXKh6oiJWlHhm+o+YV+
WJR6FA+4xvpTqvAA+/24yAWEIqHvvQO8H4T8SeuswfrX9DgnMkIrJq5/C7mEje5xav/Qbdp6wr8c
n1+6nNiYC6Ly+ktIEqGrDdfEbMGcOg+rdbFrlj1VFL7DLN7le9aKO4S9GPN8kmyhIarx8N6/msb2
CBVe0tTUQ7D1xZW4IXi1lvhgudcYGcET9FuWIpajVw013WsrLyfNIfvFARyjKFJ6GqIqA1UMzCJs
K7T1FFi/08dpYbX1eisloKX4FDacWCCvSjofKweZ3qYH7OrK1R7ofzCxsJ8AA1qLXBAwbMafm3sc
/qtgZOTPQ0PS5xNQ0s2b7Xr3/iCBfyyKY1OblE1madVJtoanbe1kL1mf/MJs0Kv6jqkTrF4lsc6b
X8JOQgYkToTWVI2UNBZTafR94i2JoVWxb99klN5fz0Ww5i20AqMiwjp2OqcsKKpELGDA5j+45ebK
MOUhdlMdA4fasOtRODv6k2c4zPhXjy91yMWx1Ik7XZdWmAbI2mSuuDrRwoIxBPbykNMJzUZ6lm2o
/9LZTjrF8+tmxTBBAxMaQFJwLJH7IJW515eW7SURB1BOHM3A9UFxcPqMM1MgVOF5QS+D1rVvRHHL
44LhFrNrb0njzo7cCyBTlJQ5PVVB7GswhX1AeGj3YDsrKz3/RvumsiZxHWC9ywcb7jikfpPTkdSu
Hx6f2sXYNZok6ChC3Y/K969A8p5xKtfaIAiKIOeRe+68/BWjkZxiJkcWexg9+A4vw/qa3x5paEp3
Fi3j9Wuti+7qAZ7fXtGcknz1cuGRClp+E64tCxpnErQbMX6U4sYADCSG3TU07lKq7/pRAd33qFhT
NUu7BCgPCl6ZTMWiVD1wXdVZHjbsVJXJV6Y3KBJvXE3yjPFQ30uBjkFzsON2BUZEN11IxUaExqe9
OvksF1YEbt4UfiGw4qJ3EUyA6p/PUMAOAFNY5QldGQj7308UVw0kh6/mfn6qV/1Omg9UvPsSwDjE
rRqJgX/YR1a1A8bmYJcXKy15i5o/l3kwfa63SnQIyRhM7RnMIOdIvNnrWRW6s167Zj77cmFaQEDy
r7pViiHaKlJJsseFiuL5fWLPn8eVpEwzZa4dQwdf2IArUub/EojJ78k7zM94avknvwothX6mGbAl
AvW0Fg3yb1F3z4jokFHy/uXqZ0hCuhhR3zIPw2DG25D48VFjVB6vFlOkwBbvt8U1ECPlIKkKEgUf
6lgTwtAYxfn75aPaJYZr1SrTwGfhBuRUUoF+vBRgqua+GYu98UGiseRHVH58xs06Bwr3JDBSJd8Q
B5f85LntkRFyeh2t5PPjFnYxtFp64BvifiVMZG0zjenyt8wZXYjnCxXxnoLTl9Ay3dxPsBRB2c0q
ImwwAdRW91alzHWyofnZkhWJz/MH7ctIn+U/zt1y5YLw67wko9n1Lxjd53QClYpwjVbog0d+dWTK
ZyVSR8PphGkz1GVX3EYpcu3uNgteZId2Fv5JMALj2PkokqWSv6+2e320lgZn3GXLG9JB+r2XUgQC
KitwksH/YnJALDkSXQR8c73oFQFN7QZa0JOZkIhCzrp/aUhcIKrGlugujJeqYKHPqEAHnl2/xg3C
nfKSqqyH4Tuex7jRLw8Gr+hqufV+uxG3iAb8/McV+b3YoG9enMyAD3tNnulu43y4CrbzOGBVCABr
LHSnsOxbH6JN/zBg7LoQVSw8D93pM1CC6A7ld6bUA8W0lHwgfLGm46Og1kZmyYRVXuV6QPUuyjqg
7w4gekEptQ4fUNVHPMOVcpJd7I3LMlwkIyRJoyhJT0XQ4BRX89phl1Q/Pf8jt4o8Kw3KdEJxjNUh
kG0ZfhHxrvWJXO0KEjHAV3I8MupVDzKygPtjxzRQ0TRUeugoE3BfTVTKzc7gMRgLoqklRbXYmMQA
C2eH2dSkYWfdDlroz+55NMDSkXzilhvfd24tZjXyO74MP208EINzJ1K3h0TfmZ0OavYpZskmrZND
N6L9iTuEehTfxfNsMKtFAA4VMMr2+/Gs63IrkG+M8b6ftdEytjnCSOi2T/GqLlLFKF+5wuAuJAc7
OuqZWlcoWeGFh8YmPwAjkz+Cor61ji2G2GbTJGPfB1A8hjt0vsCMNsdy6NX9rDy0oJCNOpi4Wsxj
sRKvLspFAvL840tFlRz3d22p7q4rZ8wVMiC3vgz2JnH8Awvk+CIjHphM4YPkZGo9Uu1WL5R2qafv
HG+JuFJNvuBvXZKI+VxqSkt4ZYmijkLuMsD08KVnlEJ3TSJL6yTma7D3HBux8ZGa/Q6oUzQnEjpo
boyBUbH8yOvsCaESP8tg3HmrjZPQaESrUTq3ss+OT4VsrYzKgjW3PB54Fw3+knkbaT1gPTt2wO0R
YuHf3Pd0MuzR61fFHOEKWACRzkO3PZcy+VFke2DacptBQRCDOpVLC55fNhTdaFi8o7nJG20GK6Mm
pbuQip0485wYnXisftKnAFQt3/C19qYEGzI+CX08aVP7zY47NBjIVYg0RLH73/hlwHt4JMJ6Y+PP
ZfO5DDMlbBfeM2Y4+788Di2rZV4zAjyKikfi138144erI1IBq+Dp23fuHIOlJIRaqf69kBCjy9Dj
Wxouonw45D1M5e5FKgzg3WgC6fWk7TI1003n9FmKHUqoAdJ7oolily85ord+Av50B5akKKZUn+d8
avv6ojFG7P1DYwzLPHmfUz1pdC+uBQPFWrDF1mNCYZ+QfhSps29jULJFs0M5tWNBAGPe1an80gCZ
Wk0kO64wC2CT1Tddc/uxigQFJGgiRKLzBHEb27npHN3fYCXwmCTYaTqsdv1Si9KdGl3Rm1lFQSut
JGhxWX3tkjNew71P2m/Ww9BnMY3aYDV+ZjSLqxAMDPBGluu3B9GiYCYzIBN6fImAtKaiBl/nE6PP
ePCre9xQCDC+hnMmYu1BaMIqH6YyXtiBlRAOfCigR/J6lXCsbQK7CrudZeoXmjJkvQfyN+0MNlKF
bWO6nE1BxFmMWaTqEfB95v6u292D2wd6VulkkCJZ15jg7Ij2ezMwX5d1xZob4aFICC3j6yDQS+lS
EmKVb0zksT6WRTlBkbAU9IQiGkY4w25P5sSvj7K/rfrzGd66nvKkYptekfABLLzAVS1hTMyiMy50
dxqA+goroXEjU0NjXBtKhsT38vo/JLCM2EWpCxWubObNWNJsjo4oi1EVBzcggvmAVBNihDKYPvqa
yjDCDtZGx9028W8G8JMMHcBZETfYJFnTIBEnFKPtyvRzyYbkZMV+fm28QtOpLu6o6YcH5SHGExNH
ncMUPeprcYjr6+eS7DdqrG1xoatCdoKh0g3/c5c9NP9+xqMyI4WWXhhg/k4z0iPoRg1fnqN49EOR
uEVdRLvl9lHSZNZ6f3Kl+jW4LyYDiuyR7Ey1TGhLIwbOh/ow7gG5vd8qGail2aj6ZRN2KrZ1y/dl
A1j2UlveG0UuWi5g//+OQ9xsxdFACUtnuyITiT/wZAFN5GnAiM2V/bYrW/UqYY4I8vFg9TZ6aNgf
HaUswiFLQLQsb4kW/Az9jbFLWMucEPSa0d5pQXoVHxJNXAwzLOm80BkZqaBWw9BCxWgngMTQ3hR5
tF3tZti5PGQoysseKYfD76I/scTWVzX871uDjeR2URzhXWC9F4F67H2YjM24OLsgpsFBoRiq1hly
wd7RLJRyUB3LBNgafkkCxMHUAyfvOdTt/Yeou5o0iKiR9kpeL52KbMAOXbNXETwTeiXwzBNicBnP
FHXJClOb2Zm07to6gPnJu7bTAcDaPuqGVzAzLmvhlqkd6aS6ODQtIyECIVgvZu0Jrx5XbYig5S/L
LN5360ZSWuPC/Z67p44awUduzs/CeaNQb5ceynEHJ3BKzO6buB94xsXVL5ySBoOyN9lv6PbMx8SD
IBdRqy5NbcC0ftgA08xhUwN5BXMHu0STERh5zHxYOlgHzx7jOWxDyy4kTKLxAaj3lOTDpY6gkkOo
6GZ93oaLccEXSPUEK0CbyhIdQonlxapX3YGjsnJarBL/eSLof+d0VnkZA3hDMmn50ntVjlL0Zz9Q
TgqqQFJMzm7kbvr4jD1tB4UtKZ9oNFe8CuMq86+5NmpCBbeMPEHG2dgeY8xfM8DxexJ3Ysr81Ib+
MeOFMZtFoAhVvEXiYn6vHTlcro7cpw9BaXjcDCAZ+J3/uZpdTUI5zZf3dxbCPBkrDp6GjGNGYRg9
dIgiLXHcJtSsF341a+fsLuUQI3YYql84IkxPWxd14ITjr3AbOBk3hLjWKBHWM0Fu5eoHVT6mPJNm
T25DSzoLnGqX1I1ZTjpYs67oV4UVl057BGhX52+9ku6WzjwuIU4EZ+fgR3ynZgkOI9R/UgOW8IYQ
ePbs9TzylbEJvBH0bkaXQDdTZZ2HcPvvzlmLz8AAPDyu9eVRkPSVyQeH01eUuXRXUX2e3nUQWOF0
dcJpm5H4A15Ptx7jvFIxOnDFtrHQkBJVPDuiCVBZXYpdqzoaqg9RRbte7/B4ADkaC0ieUlF2z6k3
7r2RgHugsuyYA7zpRUlyloc61xtK0SppWRNm1wHLaYddSS7I/SV4HKab+b27UsVJd8sLSh2qL4CG
rK+4qc/qd3vg3qvevfvNxQ5yujE//H1hQUX9HgCO4MRI7iHldYyAay9lbiT698zRrZcIa7F/qxeb
qzCukHwfHJ2PgqQa2s0AsZLfEU4cTDvDe4Ys7SFDXNW/Y9hsNpFs3Kf50k6abFnJ3tviO7W6gcqJ
aA7Zf2SPWsg2JgvQ4X34GTmtJvhGRRIxC4im5G2BMBlFvayxMLP1nGyL9ptEMIiK9eUvaiIfArHI
uyTclhDhAow9tO48R/Q0i/pFLWMj2es6eauAaKBaNgof20kYvPRwRYnRuG5TZWzbgLR7cTckfbH4
ESmMBNU6e/QA/RKvuYXCdOMm70i0atVT8kqEC1cEDz9hLiqCtAIKmWiW8JDZBcum+ZFkUqe6wkaH
cDbzPFSEpga3hUn+TWJwWRFITFFFN2gYRcjQyf1wgVhq+UWppQjw05IR91nSoyMEazY/f/lNpos0
QajeZKRLJGNrUOdMbgCD08SE08/LlHQ0nJ7HYpfaZSDSH+wj4wcou5qiRpd2GngYB1BYrS0nlTd0
4f2iLzjhrEH4Y91LwFeURCwsDI3cdBhlI/+OxcHL95VNpgfAfPm8IbUdWt3otN5V7ZT+Tq9bJpjs
/tIMVfM5t2Jj3+Nw7Y2Li7LQ8LMdxohqSh6AFkM8EjgVevR5Do6AbOS/iueJOsZpIxEW8SLJfOnC
Szk9O6BDf3qPJu3r8Z28wcx5XredZSKlMVIq3de70H1b03zBdwhnrJ1ugvyKbSfekA9q4gJ/fqfA
rFBR3WXWdMSvneX3dTTG6qCjzfF4h1OH51ZR/I1Np0flFzF1SifRH2eFg07mbvG2QRm7LP+YNzi0
fypIVn60BOc5treb2TsyTyzp84T3vyCBbURBp+u8fg+geBFk3vqokTFD6cbKkZ3qbh/IOmv5LXJY
QTkpMGMIeFqCGuyenlZbtoAj/sDfKkbUC/2QZ6fc6lZHBaJC2gu0yUzq9Njtm/073eHK87++7a5u
Vtz20PG2f9FM/X/I4d0uvOVpjgkalhtr0+wcGokUFq0BpjBO+tFBT9lYwlWsfagdVMsAu6OW5fCW
rSFFyMG7pDc27pArtLLX39hbDASDDj7r13BGHphlSbW65noRyz7sXNZujPtxOpCGIskmRge2a9vk
l39jjd7+SZ91dqEv9GAF/RNZokogYwlvmauI6IqsTus3hLFYe+uRVJwfOQYJlOVJYoPlRTPCBcSP
Ckv9zxE8ZUYvcPCblNTJfWDhgJOSVh9sDyS2WUssRGrs3YfYBLQPVEYl8iXK2UC2sIHNo6zFUqOx
tDt4+mYzG1okX7W1p8y4n85jZJulKbcQHp+jphnYKwT17nyYBORbejI6A4LQeXuoZ8Ub5fKxOwNx
Pbih71npZgtqCwfgjFgO3gGsgjM/cYPC05gWYf6PIwTROvnbKL8LpYdKW8/AxlKeMiIi6CmCOZCb
HSBwPOtoRJx5RPMwQ7f1Lp6wha9eLpPSTUc/DO1E5stXBx4/mT4pDAimstXUxZPcZiq2lvG5QSoz
T8lYdHFf0gaK3GCNpk7wgEenV1rfq59MnG7dxzR4w/WDeQMUHsxa3zYD9iBx/bKola3LRzy4891i
y4M6MES+ZCW7lCk0m5ukzI4L4N9UjXxjSv6iLkSBPk8At/rmA+Gf8XqMV60C0s9UKSahWgqs1XG9
lfWtTBt+AecBTowi7ittx4aIhXZL2uFSSchkMaF8agGgsA4yeKDMURPe023lbG8x32S6HzXIJUSr
CynZ9LZBdkJ4TWaFUI8KusC9nMEsscoY93R43FV0Z7qAr0aAdZzQLRIa/KXAyRC1tC0F0J+VH9uy
OWc4wr1xBk8WWglzHB1odil2sjVNcZH5HJmuQygHQc30jD1DLVEXLZ6hLfuVSzTPKVOcOyX1RdUV
Uu7bJShntB0AYZX2qDWF4bb/cwpJ+7BDHrOkiFo5UNAqSzxDGQx1Zwlq/EPEvS6KN/0idoFYOAB8
BsfUWAKWSE9YIoNIn/vlRGxycdd9EQmUgaLXY+f+eq+Mb3ny6txRYbKn4zmBreWeW60f0B+W25Ui
1bE42nLPFqndz/G9MKufw4gaPEStIVI0FOJHq/zSGbVp1nfInf2Wmm/1pZpc3qQjepxwUOCXHpaf
y/NzgJ+VScQYBd5Y00kGLHwzop65cHcd68+s122qDf0Upc8RiLo1gaav0UJIz9aA60V6bnC9RIaO
ZnuHa9UBqEQqx+znDW5DJudkj55vNocrYGTlDGZ+XufV2wJ7zhVHFpPJeBAXKMKdi9P+bEZM1vlM
YHceJs9SKc8aJAuz/6xRTHUhp8ItXLdQDCC0YE56xpZCvYlzvUEKantixrSpRmsxS9/WdbthHBFu
7pVIDbl6B5G+PmkM6vNRLhCTtYqd+yl4grmmZRpQNVd9veIMSmDvnQVUXF3opE+XlnAt/jQnBFB5
aX3QX2KGFQ4fOu0C51jxFAHKTkSO7o6nRXVJnltSh1eMdmDgBsYMyLxTHBjInu75fNLi4t27XuAf
s2ZSevtf37nwM3YY32zIIoD5NM95+XbzR1DTZM9uxyou4+tzW/Q+oqetnDXrTRM8fXn6AIl29Fyh
axpHncch5eidG+oni/ov37Ql/2oI5E9s6QJaCsn8QtgrJsUeEVbxhI1KvoPfp5xpVImbTpHuLHUB
LclG5BN1D0EW+lSZPw6+wmE4wSTrAUthnxppgtXGFK9eUf4I/Rk5gp5UldClghgYo38n7+FIoj2B
zPDsj1WRSn3S8W7uTDS5r84Zk5Kiuin5mSp/sNCQoNWnrKXNuT8256BjpwLg6qr4bo1W5vrskOr2
8Blkrta4ZIo0zGhLVUnxk0YbVqm+zf83ZiRQmVW74SEB9IffZ0PmGo8Bi7bcjpHHxDUehRthiVLu
T9tHOitoxQv4eBfE0EhQ+NsvDgRx5zJ3RCcHIX3z85xDj/NnwNUpZp4+gZ3Q2wxyycTJ8nMaMQNg
PpNsUqGROtdwB0eM/x9j7psd0Wa0fixWuEIlPrkdSrROR/Fp/wDYrwXMQ45gQJWq6ECRRho6FTP7
PpiXbFYPP64T0n6n6A05lvfIo85p6sSGlWMy1jajXMHTPD35+ZjgztDnbvx86N73oiDzMb9N7yd4
9VQVXdDzWd8J1dZcUNfRTcqGmYbSzRK2SnHQycgPzGj2dNl7QU1BhE9RuF3IhoLxao9bESjaeR5v
0BHWZZlzSrgQiYXXs8mYiI4OkyXO2YP/DUfGLWKWtkv5pEnvz/In7A93a19nhgIUd72JUAbzcOpQ
j890gZIRswvW2ppkQBDfhF2tuf1iqcLEr8I8HnbE9t7jKyFsf6caDkuiYlLzGfXS4D89vXqmM3fM
JV6rC0dT0ydABVGjhua7LqI7LnCrnw2lltSvNvJTTS+/F9qkK4lCFxiY5PkBdznbAS6orRwt2GlU
LK9TVCvWcAZ9RW4SEGLWzKO0gbyb4SRf+yT6I1WlFqjecYLHmyq32NLc5fodAHbp7KhgvhiXRplb
YOPj72gulbjGTmpipr8pWfMt5/XlctTbwlwWre3IC2ahBGTBdS1vipcOHsScqSAJJltoYlJENRgx
OftYRUvITtyTMbJponteVIek8dzUKfA2wyEGXaEEO2onRae5cyKxSBBNdB4mPt9iatCB4h/5CLe9
6UvRVfi4Fd6GfDosxqqgWiPxJ/XBSzgPu871WXs5TEY8It0bFn9xDv63HIMKYtWA6CcKw/XmqEzc
s5L2pbn86huHneZC3Gx02m8GxZjfAbR8+sDAXWZahp6BQZNAIYGbv5JYR4FQjoZvol3t0t977Nv5
dp29L+mnaLrGgATrA4qmp09I14J375M3QkB3lX8Y4PuNFf9lMnJbJN5PIGxdpMwygsNiWufq5xkK
XsM5U6jVSDR3mnFAG6+p4M2QpMkCjt8sCChxgOBAm7rhkl6cM1cuop1GWc7h27hRCcJCabIlk41K
MXTuBvI4DcKkX4WkYCOHl/wX7xZUH1numPbgFLndlj/t6NcgyERKF+TOr4EK0VtmdtAKK7A80vHi
J7YH+uaamS5BIS8ePBuuv77DfzAEXTuZrKyGGU/mf1piGfeY6sbGYPfPMba3TdcEoKrPOTEXKwtM
lKyY3qWev9OAvklAYODA9SKJ74Y4BexuDi2tAfwgf+jaXnc2nPTiaTcplvAImKKMbwCClUDu8se5
PdcJf8iE2hEBgBzKD4OumCusqLueJHqy35CsvdLVteLWs6+3Yc3krpypNxPw0AIpeTFxJA2ySRSU
o7oWBExKBvCV+TLGKoHmRxHGv0jWAJfbRC+wjre3FZZzIybgQ6wq/JNnWB6LbVfClBtPQnuxySc1
nZKu31tvaqfyz8NS8q7b9CQZbiYaYA6hw8fcqCNa17PTyg4N1l+7xyDyvIAtVK76tuk3osBywE8J
/uoNLjbVspXVkS2sjqx49E8BqsEwrrY19Vt0cnNBcEuvzRuq2Ecmk2b3M1uWJdEORYNaCfgspTBR
QQaCXfoYZ1knLUHYrYEmhxmtI8o/YxehQ52mBk0QhxLMJxFXT1gOyObQlP6/ORMTNUZ2C+0rO1wu
JjAKnCIgKn9kOFtd4fRhnKgWOPuyHnm4GwOuS6WbAH0lYkaENLYkET1guiq2Qdt4o3la+5acUac5
cBxnQShRM3syYwiBV7eHd0GcL8Fk3XGHzYKpv7DQn9/fS3AWxo85Ph3ZDkrg8mA2B/q+M14/K/fT
ymKF4bJDafCRS9JDchMCjm6HFsc9LK827hV+x9ZXb5c+9iWBU3LMBLWcmg1CRDgA3zVjKJUUXi4X
/hOCCuwe8dax1Oi1pk39Fl10QlCamyiN6JtKl6+XOdO23jtIl7AynvuFMwAxP5YdgBlDKRBwlX4l
g5gGBN8A0VrUe9rPlLJV+YY2qhesVNhSWPr3UhzVP3if6cV2EgFhDcGP1hufjeuUj7GzUw05QpSw
AnmvlTUyWO6qpkpyI9x6VU1rFiP0mx72zl1oM3Fn/gz8FeDbE9AIRYWOgPu8a+zf2gVgiCOpTR9q
1O6F2k1g4Xtuxsal9m4IkKkbN+GRqhmoMpbHkigo75/xtI4upkru6TV/2ZnL2+1UWTEuHKELYPcb
n/H8kzlCTP3CSiHXtR1I49UjqOhgvigMzIj5J6Mqvq4cUPMjRUSbceT1ftX1s9dHAj9WjMQ+2gtM
EdTpGOmph7vwB8HVB0ie9ufCvLkBOo/1AGXK+9ovfeB39wiFUHOmpCGsZNiIxDHcqx5qnj1KSdo3
UwTJXKUwAAkkhz7/zyGjYcN2ILLn6CD5ja6P02Dw7VCVXOWWkXX3f5PrdoSsSw1mdxM21r3Uh55o
O7azZlq979PXSeo9fLZJzkcezSQcJzzUpF2PVRW9Km3MWhPiZ69iGTlFDAx4QzXG/icguD2yjGaM
/jwdk/vqlhIJxEpdCt0wNuPUzUiADA2Mib8VmqIe09NmD376QOnZaXK7ZpU+TY2AnUy/UZiAQdhv
9DUkdQ7KR3vYwulmwXGxZK1F/ioMgVSdjsckfuEcmEPA50MWUSNeiy1cRmL5Fobu5XNUHfjXY6lo
bB4jqrfiJe7dZtyldn6176r5Us59P0Qr2Gi9WvH7r1PhvWug/ICj5hIf7MjH50iSWwiFP73+0nlJ
yk6pJzP3CQzp5G9bPnm1vfLrxHRMnwBrVEItkQc4VtCP7iFnmu/3UwVuG4M+IGn+PkynWQwXbaUF
RxMv4lznYkBF/g/GVa6v2TRa6rAYQOA2xP1NGSLm8wKgq1Ar/IQboXBQwxk4W5dLmhBGaCPglQU9
XBqDykBFPKBTRj+DGjuwqaojU06bFK59nA9tMEjxvlXfuk7AUkq0LNFd1KZJwF8HgQhLFaWqbnZe
i7rEYfER5OToNOgBnminXwr3qtESWNz0MzHayGDuGbi78QPNyu2c/Rk5nNWUEmk4sXopqIMP6Amj
YJVE0uUBMRaas51rVQIexiYkkMMrSc6YCYNJgJ0hhXQ4bjEmQYH+sdNDIXPYbnGMbp47td5lob4Q
w/OKTgp0FlPlrHk3kcH10G8L/0rR8i/p6TJ2yiHfnt6tzDrYMEhyV/cmxtbujl/zNiuyyqlsFoQ5
v6/gyZqm6TP2zoHVWDhg4y9AZYeI0qip3sGOCaGZptbif+kgtDKut4ZZvHLZfM6ZWolgXnQo/pXZ
N3cfQlQgFRMNikENY/30jJHy/5CDX3Uqo/5JqqcvmpxDHb1iaF5nYHk2Bujk7P9ZWEtUJCC3+/0+
BbgxS8LSG+TQJwBnVLCNaYYewFH6V/h9g+HcGfxb+7c2ShWEiU9zAj+TausAHzuQ9u3HLKMh/LJo
GUq8PTgzbmCHeF0+WZ6oQrWSM1kFh/JEwVwhEFQhuOVCylYVhsUW9PC73gbRgXh4R82IA5kkyuVK
yZOP6FJD9x8wK5h1Q58mvgHxgJxMV3hUlz7HXWQsCvculXJh3/m4Rdfr17FcL+xbVNt99x5mD5Ib
PvFxaCaayYVumMv4Ad6GSf5tipX5asoDftxgI8fKOtHMqL5nf5x/JywJXax/B64rea5v9EU61ifh
ODzGxVWDp4yV3fF5K9HHrvUkrFYgv3yp1KQgN9vUL4HZx+8EyXT59h2q/LmsnFunXrvh1IN2Rxyh
Ajj+oZVsN5TcdjNwjP992fVrVp/fzxPrziuDP/S9ARDTzipkqNi0VR8ZJ+MLzvpSnaTX/4BLYMJb
Z00x02Ab3b4ZFDvxcrc4MXVEAxxMgMHbPL+TfA3eaniNGGZmdzCBR7Xzu+2V19yMgC0uj+XxNMNd
qgAKE0Qc7i1mQoL6tQgV6HXy4HocQ63tHbNLJAzcuZm/0Ei1RuTUsc4eOll57geUZ2NbqUshUgW6
ZWeJYiAKA2i6oROFuIf7YeEkrw+aNSSWYW1Zk8wqds3ieGiXx6YA0+gI8WFxBSRbKBTAoZ7/X43U
l51jJUJvDKV9b5L58reL6sYCQfzCgZVlsAcR6ClUq+mZ6UhR7R13gMdBuiu9g9NLup3o4Thyatzb
Pt1jAlXPS3eJYQGEyYbMWjysy6Q9aF9l7zmSaf+c5Nlo1oXezvIFJnTPjb1a6R+zUqQrd/DCfTDC
zo1Sx8IVxlGqZC2dSdsNCQYGK5pSB6TCGrW1+vsi0wM9PA4nsgQZG0Oe8zdfFZyTkuTNn9rgd0CR
QMYYqLhZGWH9ba+VSJhM2qfLglsDye2tL4Ss7SGA4b0VMN3o8FcgoUtsJk6qHmv+0ltJcHb5mzrm
6q42rOtup5R647hw7ZDRcOxXBZceQ3ApiUCvCiLLHQnCYDYLdGJVQT0OrqBEmpnBcw6qqFcTOb5u
nDElptEcuRfYIUD/wDVFNTyRBLFKfHATEFamLZyODWAECgbv3OV2wdz1qSxb3pBbR4HBljToUhXJ
0Oee5IjB1uHXLvqQsrQNuIHUpwRPiwPgqTlvsxk73SwrT2+4fdpbgdtGjoWuGyUcdhpagFTt0pfZ
yvOSWCnvKt8iE8KkjMseI69I99qjMIVEF0K6z5lG7e+iw0I89Ha3dv5LzHW3s1vnyk2LMFqx7dLZ
Lj8GDqSUcHB2nT1cTwklFmiQp/0URihU3T7RqpvipeF+BLceJDkyHFL1cb4FWBEnjDp7//06Dwbb
dTl369phGTCmHGwuAfcCFTYPPqxRah/HlF1Eq5cZv6AYDfFMP5Z/rUw66wYV0ZoSteguZ+CitT/i
pqD4LFx1TDQNGZvqRbKXtAAycZS/j4hyBX5P3gw4O4PSCFlTCyOkwl/Fpv/KpIiw/RYJbluUZCqe
f2xy5VYE0R2fLaPXwv+8Jk+gqWU7HMHSxCDTMaFBvcWPf76lN9X5bDU2xZRrPHfhEl4I2wnaf64h
KoXBCDSJrUlHrYGYDr65uSSY6r2FF/AV1vW1eZf0kqQKZax92Quftd12EVLcm5241CxwL/SSGa6k
H+HiuTKLMm+tWsRnqEkxUxeKeJK/lcGEErNdhUJnWeGSdpT3uws7wIG6+FBetJigYxI0xsnlWQ+b
O28amh44VJ5yVI2mxZFM+kGVCZ2mxGhKeQxtYJzEQA9EywByH+QNw4BjgaaawSzh8kOsO9pQDmbQ
JcEkQo19AEbjh3HkMb9RPyzgw3eoKDyAyzFSGEF93kQhcfR4UBu1ayRCPlYsLCzrkmwzXQqsgtod
DHlICasccmYZDzJ3e18FydB/LhZLM5ZfvbSqUb0je9c6f/qCJ5hmEfZ8/j5KwF1dyTfIZBG/KeiC
j1sOKzHoeJQD5rntDNKjHlVM5KrZ9I7zJRYMuShUySaYyKkaSQOhyEg8kgFkUGGgwG2gI4Z9e43o
94sSVRA2c2P4/XwqfdPjT34aaP9hw08HeZcYE9QyT5RBZCT19uzairpmW6is+Bb9Mmf5M7Ja96wz
wufwM6zvmsyPNg9xLsUM5PXjJQ2XJzCrYPNm6t+Ogsi4TS2i2Us9BIrZwdg9loOkOSdS/bc1W5SB
B6LJVHaK65AAQFvFxbxMUJgzG7cE4dwNsqZsGEgJCYek7NDw5wq8Mc/0hzmAE0oCPG8PIcbGKE6y
gAqZvxB2WL3DQII2BgJ7zeX8r5qTkGhu9NFWW3gBx2N+NdZwABA1xQuC9UuHRmrLJ4YlmSuI18MU
VVOiC3dBKUOiNMeUocUoB3sqSF9uMcDm/Rd2KYIwmdAFAqfZ9DWXt2cmh3td6t3rGVdhan+v1RO4
8SvaJl/lE/K6SOHFJI7dCWdZjV8hR5QVwkXqx4IkGDbcR4duast4v/GFx5anllJy8czpfKtemr/v
z/MpwaOQ+A0OUcGnlJMEy3wckDb8tZr3IDB2hh1TeM9JPPwV5p7zvsCDrWKDtkYXorQxoP0riwFz
5yn5w/s1RScvg7PxahpKpitv5Y/bQ/hlCs8/ZXbN8ho2XjdujPZ0L5XHNZl9GddOvNyFcLLCnqP6
ESwgGNh92th0PAYwoJe1G5oj9B5CT5ZMQT2NddvtBLgupFht0beVNzjeqMMdnxBTGvN/2meId4F6
UOlo4DAympubnNUi8ee+XDcoZewwIZqYGxkBL5xGhpfkoC5nP0aTRDowECiKgwMUTuwxPZBev+sQ
kWtvBDSl4ME0UxRg2l+uW0tsUGlmZV2mO+B0Z914RRHB6rBzJxVO7FRJuzil2TfrYLpUzWhumfjH
R6/TO2AhcaUXl1cOZssa63p4swEDOkVIl76AJDmssjYn4j7tdUO2BGDnTB2oq8t3WDevNw6NkDQq
01xjSUC89eGo+kqwlPxJ8DrlEJqv+ONcm+sjVxUqUzFhDgxo2I52ATP4Lz3AcDOmourPL+wojImP
h+5W59ao+22s7MBQIZ/GjwsllYeOAngxA8MR1NY73x+R99aTxCtW3z3fn0WWhi3U8MRHk0S4yTKs
BMX0WUiwS9062iVf9xQQ/CXqAlpTvaYlvqzw6yLwApuDsLWSjc4hReid/WeOJV46qMm6nnSvJ1vV
KhNm7Rj6tREj7lajN8jb4W21dYodZLjE5klrH6EhsGt2wlrJ9IB+BtGTG3r+hOp/B/j+90NbPduO
MJe4O1UOAiQc4nNNJFiS/UeRZS0lwwr6UA5hXrrA1LrdAM2ocpPmniChAw14g/pDnGOYmWm0P99v
OJudi6RQCwVxKRbPI2xwJ9MBNCgWoWIr0Ns57qJkvIBiYFvEWJhxUkQhimc01ASyuWEEKlwmmJVx
OxcrTj7yvI5jO5/9dixjf6q3kAdMAKCPO32jIillYDOR9D1DoZ8U9chDCxuvWlTmDLXalVv3BcNa
9GLGUv+o0q791xuquaw/gMZwtjgqOlbUUvZr+XYPxFmNcg4za0QSCQurfgTAMCrKiz6OFSXlj484
I6lgpLLd+0aTW60En9CpIWObhCI5bqDYbrVegA3FbG9J9UvmqbhF5NR9kgxY34kCBb0YuyKdh8fG
9FUUeMdga9XKGJL3Sh/hPfkKG0jJyvBTqxivfAem7IcCYfIIaTSrhm/39KL8PszgX7FSsPrXjy7i
qDwDqr3AkRs8M5OCrGUMtZFIs1XI6lxzSTyeR8eIYc9KLCMy1tgcYpn7TLibNCwdrcl1mMIWwV96
RhT/KveYdqth0mVv4l/z46Jandezbz4RQF1srHuPEZ7kg9dJM6R/G1NhJTb56zMcHx6H76baA7iP
1HF4nEben6Tf9Z8iDpxCNjskz5bEjZVaKwgUtHWlyl5XOTwXvptUzfwtz1A4a6tReciEE7IZnHQE
dVRTDlFyHITzY+QC/saTy7M3HfIv3WMOQt1O2x4dhnJ65Ww3WlC51uCatubEgRHCAg7oU0wzwJUz
t58dKlavOIgotnzZtxf0CQ+C23Y7OihLqm0z2uWQv/BUXYq/Gc24mJxwXeflzM8i/QdzZUIWGl6o
2N93cjbcGKLrAPDRCMeGCpLKxH2oJjbOBtxLzGHj6t4iml6PhR/L0mAoqZzF52Zfo+Rz+mM+kNVQ
oltpx1ndKLxli9Pmn6zB6w64y/MjUZ2ql7bfoO/AfnCSIHT0QB+mxfRm4m9So5/OBSmEFtOErZR0
kx3oCiLZt1FS3rFwFr4gMbKR0+Hs8CybCL1s6kyFf/wblQ0JCjoGGk9ip01qSofCybYf2/GzidHn
Sxq9Y140ZBns+9GlwlT1NpD3Q/1kyGlbLKJ4JkRu0zSBLvuOZBTPpDi2c+nEN2d3HHyWHQ5xh0CQ
R0Z2jh6u02+ji9OkxLy40h9MrdkKSLF3QbBL+L4fHlSD7dkhsj2WSphtA2tEZHOKMttEiZmO68IW
l+eHQy/a7IyRIe6wd9CaCGIhMfuJuU2yTZOgugujryzM7p051C1LNbArQXZL8iZCmgalLVJ/g3iN
kPCxlPl74i1hm17qO83CBPUjUzBS/VipmFCFweWgv6MSO/EZ4oOYvayqDj3Gpucd794Dl0dn68OC
Wf7tPy768gYTDbw/37zNJFGDdxSdVOn29Vo9Gn/g5ALMYB105yZWixksAo2FFZfgJSPIuG/y0g1z
VyrS0saZYptimSDZjdI4a3wf6+uBW+MZcSxseSOcJrr+PNB2NElW+26DDgFsvHr/JTPrCf/mLPos
VXqIrRNIDx6rH/vXa6f5/bvoXqUDzE+a9qcbq1+R0MM2778PULewueVzwTAyC52viIJ6E/8C9GDD
CxBDQ744YABKOz4WMJxny/+a/t2BQnqBwuosy5rKWmc2pLY1GKZyW2ClMly71g7cohyJHNWmky+T
Dss+/QSB/6Ea7BYfLvhDO0tQ0WftFKxNgrwYYQ8ZVY0VRCZmGLyFn9QcyAFjY3V46u4kXAqhy3aB
pq49FZP7/k4cPQzRFCnYlvb0dmPq1RkAhLucYddLfr9ZpO4Fgx/13iHEvTVcw9aK+7dF6zOas6le
7KNB+GhhgHhSUqPu0xVAFbK0OYAJD2S/lZHPmGrGB/P49q5FsfQ//ktFZdt/Yw6uriUYwwPIU2ys
47V1pqAebgWMoxM6ABv0XDjRkXFuO8IAvDiibM+FEDm8cHvgyeDSbQV85hz3eQhJJiNBVgit9vAX
8kEEt2s7g44yoL93LCf1NdkwFjQO/IXTNWMRE4ZQTPGHqTlBkVIuTk8GwGevU+6R+gGXbCxOaZLV
1/Le5XmFbkieCXbcDBl1PfJwxkxN2YjnCKDuDrV4P3DG8Pv6SKEGy5Sszq4bQh2xTbmXQDbuctoR
bxGWPhhh1YkU0kifkpQ89WcQi/L8X1xHptFupGZNmN9fgaw9Cy843+QxCz619Rof/IfSzd4Dm7gT
IpQUoNCa2C211kfWdhaWFG+e/B8JctqY5EqUhaexP9b3zwJveRdgzbwHPpobhZLAJrET/+4OxrGv
cKlyUHRAbFA79HK0bjNc13AwK/4N+im7HgbCsrEsqiLii5WDCAd24ydKiOiSAtA3dWegThTonZt+
DKfKy/qhasDaaiicHLqCJFMTtmDelvtmMq7295bY8q8Izlp91TyZHc8PmNUBVeJ0wn1Xkni6zG3u
ewWFZdTMsP/4fz9u5NW78lt2G4gGXAirnFPik/F/DCJtCaMSgnYkg/WCrlJwSYEJNBBt5s31QSeH
2KkfUkTroM19NRk9OHAQt37gUcpkPZ3dY6T0qEFVRcWVBEE8Isk3eLCp5dG5nPGzZ90UUT+zwmV3
HAcPd+sjbik917UF4xA9PlUxe3HZqCKoyAx9VtTbTDPl8FwdeX6RASL5mbYzWLJtRAkHS65wdvNX
xiZBD8+dWhBXbLwSgjNrDr0458FPW9DpI5VHWh+Zqiim6qjtcZRSKxxCIcesREf0BK+gdm5xlK7t
ZaengSZN3ku/O59+iZjRRb28MEQbEFt8PdUmSIM4hFaOD9DUHdSx+2hCWKDFtZU3wbt+AREEFDQq
ZScQt9xf/+QBMxCA+0fsH8WHG31GEmOkaFkeLQ5ovisSDvOHCtQkMhFX+Q/8P21pa+dPbkhhtRnz
RRKJfFtyJbjvRpfDgCRYn1egCkFwYLbd1XGkPnsNELj2ygQsgO0H7hKKorcMVW48v6ME5nhr4vAY
LMU68V977ZENctjYDgoxZ/mR8ft6ct1SUesAUHv4ABFmSvm+5U8nmoXfz5CZre3hKuyhw1qqW3Xz
h08sXb7kw1GbrMuBaZN2ZwGlwL5XR/fnOCLMCPI+lgDRvlAKHoDwQiDSleNr9EDvRdsJ9BX7D315
isbTOGYhFCVSJZEw5ISpWm7b2RIqk51CUCvblfvFgKHvoLJqRFg4P9M69cf6Vl9L15/xRtgcHzBy
4S3syqTx056WDR8XtjdriGrd95GehgrznuXKIw0FaScnL8qzXelXyT242LTAmUYIejwq8Eljseha
oGloYYILaLft1PqmO84c5y/hNrTSBYr8vlWGy1ET/mfNn0X7YidBUklKm4wduPpDd81E2wTADyVx
7mpVaBMgwPs+ES6QH2oaTxvHPPOiHGz3QFFIM9XJ+UQGQ8alaVujhrt5wtxO2Xyn/MiyZqAUe4nv
y+amo6PSQFzRnNZP61wFd+15pgKdmF28e/KatEdiGkU82ovE1SzTC32HKusGuOFi+aX/aLAtELZY
8IUvnJmkk/OITGmL8lwiw6oP2nMkswUPFR/a0EejLO7O8rwVpfTSGyuOkcKot1r6etnHWzD0cGzv
bNfYMjbxbWAoUshvGZK2Oir6njIdBqwDgB2HDAFv48wB+oXnjJm+KrjwCQaEi86OP9mgZIvcTDVo
Sw0TmI28eHoNLYkP2Fk8VibSlS566Vx4AI1fAgmSs6inbhDe984H4rC/1g9CcFZ3qNxrv64g5udz
zeDNghi8mlYK2zG0+l/XhbpRcvcXnTYdr9yvOvm5hqlzGgpZfivZNvCjA+dtbsGoipJBr5stHmVP
f2JiNCoiSOsxAEgXNHyVJX5czQpKxAKdbj0NU8ZP1VIKk2YE9HfJKzm2COsRCfesb4M3qECWDPQ+
qGYCuNtwLmqPBUzba3WrzFp0qfsrC0xn+DMUME5cLdWEWDV0T72pq839T/jecD+J6rBP77TvbIr7
k6FspyADEa+IIQOLOoiFoyWPbNek6RfHuX/6i++IuiOg/70NTPphL854z1QzUeGsVPqA6zpaElXG
C1TX7RW8N9uF8/wmlFPpOujzSNWf/Eyk/9yKidcB9Avqw0vCgBuSHBkEBg1RnDChBh9nhSq0ZF6z
sWbXmyAvgTrwH+0JDivykMslaXsjsRwRdp/xjeo8hMb0U+fT3Auqe4kHwR+GWRv3zHNSJ0QH42Fh
0Wx0xdMhSz7LPMZVAAs3CUJosyMuTlf17n4B6MStax+WwCIRPc55lUjOMayKjueZz2h2B/jxTrlq
TG8ubIbMZryVOO8N2azOUNWKoC0q+pjseF40AJtV/cVBx2kBjgYjBxjmQIwJYXTI+xXaLejayXPZ
4OAikXuWFEtqRLM7OMz47298QzSCPxjh+CV8/27maF2I9p2NRQYFeQpQBfEW+qb+L1groKZxZ9Vc
2NQpcwzjZ6QM1LURpUIUvhWF6BOjYRxT67sabnVzojLQTd79EIMGlEfaQnt/GMHXEMzzs3CvQ1k1
4xnDLqtN6vixqVjtjBBm0ZjFxx40c8nJGfZYv9x1X6PBZ7i3uifdDQru+bjgSTZd+fjtElwCCK1d
Xqe+64gfB7je2uGDU/hs/G8kY8WtN13LgSSMw1BkfzoJcQb+PapNbArJskmN71BjSgqg8sv+fLUV
Eml7NuEscU9vI/haad8xdO/FTw2BuXXltGWMSBtv3bN+/UKC3JfGtK9plyMdeR0vHnaE/kEkW5tQ
V8iw/whkbFxvmEIy2uzjy9EvDKNESebbELlcIW111OxdGuRZfG1z9acvUstPhEykXccXxuVkWm9l
/aKxFviziU2tPhQbPOJcP937NuPF/YyjvIrVKVibODpxE9/vDfMS4ykX0eJf2OgBXrWaedxCbD4U
JJfHoI8/4mfS5GOj+NVNVHdwpZwmm/JdBLRkvfgsAgxmoI+aA0z243EgJqqnp3ZdDam23rcXmcZ+
KCe1k/XG392etjSoBIOK4aZU0T0yayK9slpp3iUXRkrvCYUN4URl6/rhLdtR3Du4porvuR51qSHs
DYB45vXkurrDn3HiPzUefSQOnsP7QHh6K9yAcWpc+wnhw38Q9ucrUKB2EonHtkIBns6Av6LJKCnp
4X0BTHzl0D0jCcV3SE9N/mgXcZaT/sebL3TUHWvW98NbzpueddpjDnL9CuNiKo+qatGVZQejJktJ
9U6O4sZrZOCZqNehCwCQK0A85+KOr6OJfyb3rSFt8ywfrMr6OgQZ0+M/70Shfk5vne410SSSzJBB
uhHtk+EwPtm6YUnWskSSuZsaFealUSTkcozezTyXqAGlYWW38rU1zcGH8+gxfl6F66eIMMNkCEDA
PmrAIwHkUf5pyUauYIuX6P3Ygb1ZNyVtBWTbf9BXIQUYN2u5V3gkXgYIeQAg8SyqwCeTi+ZBQSUL
NfhBRJzRBPFa7EKS5du2LmWC5BrWUYNWkhg6CXHJmsIC4mdPuClpzsoxNy24wVkHY9a1fXIIAO8h
1x/juCkLgyt/ik5Zn5UjSIEVPqWl+bFdRciwieDEa8sjK/E/0OyKePNcbHbOiMSCqnAA2zcRW0Jw
7KZ1sIkeNvy1v87aI+7Iuags/WYh6UizmRkRUz9gwUUeY1ZiiPO4v32TAPGWfWftz1CChaf40Wg3
lEIBS0DA9zERekn8oH8mGwtY0o6IGMYxrm8tbqMK11SGGW1t23rIH8dSjc9nulXGn7CUPHZ/08d9
5dUU4TM6/ode3rLv+b1MJtCKz37cxX9Y0iatkwVe5A+y0b1yAOFtw9UpfzuAeaHlFz/+oRCY/zqR
qjTcifwJx4qfJJ71PkNsaVIx2L+zssABFMI9Ao1owUMdHmyAafMpN9qvEgVo9MittyYGRm71ScQm
N8HQIq0QllaGEcul2y/vkCGlP1N9XcRVmFXlKJbtO+a7MxYPgct+jrXiWieRT5Egc4boCFQDGPXu
Gfa3182TOfPEbI8cf6fXgp1fViFIMFa90YnMrgaNU0cK3Ukna0tFhs+m2DPNgV7geBRbMyD25C/k
tPLzaWH8X1RxAuqSPJMkRS2gxgmKr3HZJTEkU5pmDl5537HFJ+iVnpKk3JYydclcW0LQE4NSq6Z3
I1BNcAMbXp6NlZG4YwPCqf68KlkmGhtvk72Zg9F4SeQ69un/Iw1DWuA11TFpYFMQQg2BvBQEbRzm
IC4Xrjhvf3g2+rYPcxgvTW1ApJk+OvIPcyLJ7Por0UO6xQbqWrcYowhY9jqempabZTTaVQFLL09+
u/huRr3v8Sl9CejNX1SqF3yvJMfqspAKJmkmIvG2cBTz4s2FYIXPSDntDiAHJpzPB8+BnCjF9HaJ
hbVU2dlR60ZZNTLorQRLevRdHrKzBGWEIVJg7aGj/nK+u8LkVeD/sQV0Ow8GJM6jpXnl4tBLOGwE
ATiMAZAbMYfra2NJSZgmir0WA21moikXaTupQWlqU2BGLz69BCyasXr/d74qZyJFWhmeNeyO/bz7
9iIVI3d3vUQjccjNiS5ovka3dNzktX9Eoa455vHmQ+BG0gJQ97mrZ6Kw3f6l/HSmjzLpU7WWTzsq
I+ZFMDhPhorXO+Zs+Ok3FAeN4e53iE53DnfUTG6QDV3PSSxDvePZEM1nl08Q9+eJgN3A0W3wdF/i
4bxyjt4ZUPipViRXEtkMMSl381tNzvxtNQPitv1PyuO9se3Sqx4EvsW8y0g0XffZlWlhpdWhmRMh
RWHR2L4qabI5LsN2a/eQAjLhJP9R/+ltnmN1Csok38csidNTr/6xgPfFy8WzzMpT196FRyHFrYu6
D1CAI/ekHZD0O1G1ZCEyUMaLjiwfL6DjQB2WNz+1ZQRZSRniuPRpxfQ9ge0Ow8vxiiZ4DYEtGSIN
g06SCLcNGjfeQRnaPUrLNLnu0PDYdNe0M53IbMhVeHJ2ZDwvFgapHqF9bFrMHbA2k7yc9tvPyB1g
ZCvJTlcCIjR4waAHOEQ/Dbo6TPHQMQAT6Q8sP2rZf1QivkcQk0s8FqMELwca3kmGTR+QHaXXh+ep
VT8IcciXliZNzeY2HPO6Qo7OTcLvFu/94Huc35Xwtnrcwqb/mO8KgIKtxCGsHyDngINbTkdYOXnR
NkjdWA3mSfS/+y1sVmErqMRJ/LEIWR4H3bOf/mz0huewDNDdVnqjWsHCv4xmDFndNuhFdfFidbyK
5PSJR07624haeTPWi5vVa9kkcCcnkfIW4EuzUj0QiAPIygPl99P9Vel70Z4VaMIg19VFCuokgJ5C
EO9Vyujsajc53HXQZIjJBJbjRudDz+lLSvPBrd1EYVppRx00mGSRjt4gi9d8wSBiOQB7LYeFmHbr
881S0p6LnO+fOmDobAYxfmufogSkGb7KBDqlojjuNZVN79GGEu7u18WzXHYWXYj35qkhFxkHrK8y
3k6mClCwuupJryYa9qQAtz0OSmeA1OPxT6NAWQfCklF+yPhLcnMrZXpRxFD1EtS7ehnhLN68NvaF
EkwY6JZYOG/0vFwRZbeiMyGjSRMOjr6wMDuidbqmn0O8swdS8tNX1vfNHdPqhVbX/Gw99iatm9iU
bveFqX6H043g02g1NHhiVoUqwL91V1m2Uz6k1z29Q6yu/EMQkbOb9nUCgL3Q9cYo4PbPkE4SaDE0
buhG8vAobYtaaikE0m2XugKHxQ4T1C8gmlnMs+pjYMS5SPFzM95aM7Ii2nrZi+CnP4dc/lvOoYEM
M8NWAO//kQaY3hQBCh5Jg0s+6/mfjv8V9DzDKbqYA+qZ2dqTnwPb7g+ZYJ6iOWCo/M+DZWcLmwpl
H2BvPckP9351HHEqOw73/ydQJJQKt9Ixlyfz3yGCl3XcIkoWhkQ31Jgkxyj7Fg+cI/EvjdHTtqAS
Uzetk86gxcWLyj+7GNBB/8Uuq96KABf7xh/rcgAltY3P5UKQGJqb4JeJT02Lmq+L09SrJh66BWtn
HHPCs/Jkg4nMnXMTMPW9+QqHZH8Z0nsbtqH9s4eEIVsfB7Lj1Tfff761mo1wfdmpUQCjLs7mWptd
7sb1P7mo2VxkNX71pbOmM63Puk36BLakCJKMNyaw1rpQi0InrV2GUMkNZjqYlqblP4v4D+1OhDhZ
wyUKM/YQYcUUNF269QLRpOgU3yGEIfD313brsqKYPBkORY+bjb5DVKdC7F8EesnNudmpnRl84+Up
6GmMDTvDLrZ05vOgjDlGRzaw1LcOK7Q4fSi/TadgBJTtaPikEfl8MMxq8E9BLOXpWDkn36YufXgM
Mj7fJlHtMyCutIa1BrBY3rF+xzhnG7IdpbTPr+focOkty26NL21ZJIBW/PywGdZ6+3p4nzZPRM+u
YKOx1g13K4opq0jVR5tgESwgy6n82IAOIq1GJ25201tXu4uvZIHK9JxhUaXbS2OQYabL0Pd1gxS7
Btc8umSH5M/N4OPF37Ah7wp/Ajojk531UXrURZNZM81vWhklZ8nSRib7SAT+6FXL1ch7Uj4fLUqC
Mm5Hbo9HbEAzayyQWoMcJnExdP+yfzxY0pbInGOegCG9jV2uwbHvuDePZSbUC8k6CfMrIskxDUOA
86fsXkpI+lGfCuDtYvNIAIRIyuB3Swifox+RHaz9rVYB9fX9Ac7D8ob9MBr7rbGqQZsymsM4uxlB
u5ZNkQnEh21pCLFSasbRQFDDabm4Z2csT6SKYf3tjjsiI/Lrqo+7poLvJX1TLY1ZZbK00Z7cgAAE
TH9SWqyK8JLjSP7bIHxn4iTcKtBKeE6i4zfNyXje1T5oWWxuXuOCfsUVrlFbGOMeU3T8Wey+DABb
kO92Pokyt1i8RSIn62xiJroibI2kAfU6dQTtIos1mrcRJlQ45+t/ychlK7wA7lz+BiWGpMCnbOhM
cZj30aznvY9+CUHN7eYE+jbujVJAnA0Tr1CpDodMWdjsHbcBkAMh5iU9wna+sej9WE9Z/ruHlvnp
SFntCB147immvszZC6QKIxVWBqL6hGJCn16//4g4o1fOCZuYb5dP+m/SMploKB4WcaU8BC8vD/qg
fCL1b1Hlcbhz9OCEDR2H05VxPO0dc2v4Meut/uy3C8u6vTXUrXE7RTqKrISC0U6t4c1koKTS9q98
qtNKu0Uut7pky5GL2IHMXHkijOIXXcLsWEk2gZ1uWqVmu+iEOIct9fYWZ1X9koqwvJHJsvPxhYzW
96X46z7TtyPhO/a5lXLZBBicpGhv1+ZcYa1j6v9kPEfWt2tjjw5zBOaWU6oCCcpMI8P5SOTPOKy0
T0pAdDKdnlC0TaaQymNPGnGAtWPcw5wBDWgiR6jCah3zZxyTAx1LX9jbS6wHPZLn5F34lrea27fl
KXwU0KmeBdlLK9FJjIOEXBRQHd0bnOmT/HbNUZI/uM9WT2xXJ8IxGknyn3dIx4QAFL1+VYrr85BQ
51zIF5+1Jz2u9E0r49Cw+qVvUPmzTYD6G/s3iwt9pCL+3OFBk7Mhh+hQ6eP+2gJVUWh3VoQ7d2Wo
6gWVjloGfQ06tCNg4HfrFhZ5Jp76DmEhv+8nppU63GLkj+FV+RJAkevjq0n1LHNJ38QAUSHQknkt
PYJFfEjsz4qwtsASBE2CrBuXhn3mhuvq04OC1UU1hOkjmKhSw7QjxwFDIA7emGrF/pVXVdxBSKir
Z9XnqaBZaMcSuSHUT1ds7sUn4adML6UDr8CENV0mZ/amz5l6QrkLA/c08z5i822sWQ4tNqzlKQu0
xDXbrSB1d02zfi8NC1bd7vOvzaf9l0eF+vGd/rpkq9RnLFnhq7htZp4gxQEa3mMSBF0kS2A4WKgo
f/UDqxB4alLvgiWPMP5H6A1DZ4oIoN3MyAQeaO1xa4lbHiZxh8W6BVnzto/Ek+WdsoVs7WQ4EaFm
xSrHsajuK3nf3f1hOhttecuqCFTDkGNZMad14uoqY4ZtKOBb2HvpufLUG2Ur8+nACpksxXAEt6YN
nkgszgQMJXOMVIKr5I1UxhxcLIfr20p+FQP/hp4hu6uT96Tway2wMvhf9onJv44mUpSc1hlFOaLS
fsGDsuR/y7MbAO8/W4KDVTTq3yLLpF+kbkWn3sDglQi/tOpEiyHSXVgs6k+7nJCcdc6zk0aJ7WiG
KzpKwyyYl1sPDmskw5nrmzAm04xdnTAWR6xCS1/nk3rOLsX4pLJFCk5WPikgBU+6gx8d0BXYwH4E
fwiZ8wx1bRR1l/wDsIGoGX1EJX0uRitikmUDd70mnPSE2m4VERy0aUm7sqxZU+QDkfugce8Wa7KI
BsIjVno50Qril2OMv8P3XL6+TBWPJ86Ijt0nBRLhNEjtBKtLR5UFyTs9otx/IDbgSr8fAGA3bvBF
PL5xe4cT8uXxsdh/m6wC+jpCwPX08CL+Qjs+O9KCLA2fKr4Ywr0y8sk1zEwugAQE3GEpH2Tn46aD
Uw1QGzkGbVyMdrPzg/nPrOxD0sdFiI41kMbUxEn1L4rR6d0wP2OnjXX7XRLMvF9xNfBxWcwd4q4i
drnBscit8Ez42eMl5VtFXRBFHUWl+xbyE+BMQ4mgLfBgVQz3Su+0bvrrM6ErFAAAOeQWn7z+i50Q
rUefMdWh4OLjMrMGZUZO3kJKB+eIiOAWSHmpNXjMccpIoHJMOe7X5vLc5Ya6ciICE4uc8+dkCBUW
MyXqCTmsl47LClcS/uLr8s/M+K88I5dy3d3RuZVXBVPX6JhJIZN+gtv7jsGJL7ZmIv7D4sOTQYAv
YQI5VTtQkeMq9rMzlOpl9zqWOyMEhRhbMcxofp99Tvudi2h1U25Yq0z+ytRM9jLSoPG1fOmq69UN
Zb09eCkDm1Y73VQ3dsxdEO/bKPbB3i1RyF/ZMlzwM8kC3ZOmoO0IeDHK/R60g96B8i3KXoBVWS/i
TwIZIFq8FjBvLrsSmmzB4Xzf98a44gxFC1uVUHD6KG4ZXRoAXBlk7LDqD2BOUBUgOyNDnzL9DJLq
3uPhbzTHy86bqy3xJ9spxikYgfM3oIJG+cM6bVclX0ZkRhN+uDEt4NBOYit8NzXj3NO1p5ZWfbuL
uo6Y0RSV4FUskDv4qyLNQHEqFkzG/aO9cWaM3LgUy95VIM3MstpIcZBoz93CLa5tk9Cyra7PaMcs
1t4ThizQmL7TIPdjdQJpZTZIzp675YisxU6o0Mk5wQlWQHHyWW5p6zeeU9ja603QnSpp2x7amo/t
XTv0fXHQqxuEuZzY051Dr0PmU9UWvXP+NrvFBkkw3gb5dPDa9fzMVaBAsvIciXAemFmSNfNV4xMe
4haEBxLgN/sAs1iuGKZvWZ/h/UO1K/JJaO68oGvArfp7SEeulCT8It3NJdRwbIHpkJV9b+WiV0hG
UZgCrWT7Ro9mtky3G0P5QiZg2UYM2GXXG7fXlpYkOb0EB4p8o1SgVv9QObTURbPA920yoeXnK0kd
LDGKcZ+o+U8nYVH127oBBp4HnPZGAB+s6mU7wBexSSzX78c5REQ6UExU7EwWVAjlX8qn1hcLbSjC
G+cXdVLzcieP5PtJhEFeIn4CknuzGbOWRE6wPYe6QxZ5JkgiQpWaPUdzCNNPGtW9EkcLIog0wcOr
yJOgptB8OQ5PTFU2XQ0Y/qFcKjrDzwR2Z93CiunXJESMylij3W4bf/zxfg4w+5Agcx6JRpOYFuEr
rKCY+f0RUm82rPFNUuTKOu9u57wKBoKsRWuh+gWKZJYtATaoucxvTKK0L/YYpHgJIK56t/MTNqzs
1iQQUo6yhI/mdRB8+6TS+qd4USdY44xPTQiZdiLNJMiXDaUa08Np72Hbhts1V70JpR/hNU9E63Dj
IQn/gm54P03za5t+M6rVkJd9rSF+vKzherJGBJCrhpuanlaKZw+kJ58rsofidjan6nNOv21rnUi7
2xmHCcsDtAEsdGgyax1iHqv1XddO9TNu8loIND7HmhLww3gbmFvbD0kLjCGpdxFgZALkKEOu7VMi
srEooEnMmwCP/1J0aLHPwAR+H5Xbs76Q8v7SPlaN3QjjTTD4s6TM1acvOMxq/bH/ReOC1kj0BDK0
VtGSpZeQAOuze2npMyvN0JBJynHSBqGk9nxpe6eQJ0aRJFJMhJh1lAIIYmqOYv5Ux7jzVkhNZKOg
b84SsUGWlFKO0/WjjUoNcPR0ziVi/vrXb8AIreOSbCV4wuR9aCKMmhhGoFrE3blpVPbwWoIei9RF
cVvKkb0YAeH4rhe2QWnzEUl/wy1h3JSbdQMBxVfrZfKGqFDZdG35O7nU6yZ7xJgsmcrNgiF1p5fT
Z9dcvukFx5T2xhvgpPzVnUKNmD2EtLO0F+0pyOzanqKSj8Th6GeyyrX0xuWXZDXTha8qtRqdjOvG
DhhKIg7ZMsGmLT6Fz3pl8fEBA5w/4yiE4tN03s4D+5LWZedJ0VomMHAvPOP+BRpgkaq6v2m7YEcy
1leQiY7YyyJqVvA4vI127+x04HVuIOmQFmQtJaSTih7X0UUADhDSuQEc1bgT6Uz5llV3OaEayiHu
QNv/28YYIWB8gXNXf9U1w15uSKUs5Gj1Shnz9Gp6B9qigeD4LUQhbreERwe9pol/eS/1B6x3pvAh
sQcSneOkLFeWMSgK9v2qwVcUeqYkZECm9Q0usL3BT1vTwduGkvoxw0qiZpkrz96PDDvDg92Tfqux
SznwS2LhQ9Yey4UiG+fyXK+bIetKcISRrJfiYAKGyjwDOiBXCpSgBXPDIWloBi0rkPuhJpcp3PrJ
qlplztCugChUQHPW6cVz4yNENpjylLzaoRAj4oNUqp6P3zrupHMUgbEeTzDYHSpV9Jf0oCBakWEv
iMZvEAaeoD487ZCoD/LKxxm+r/TZagVxrpyqpYEKiNLogkTm/W8kt/jHb+0VDcF2t6LsxT6hQZAA
Z2ZAgoM7o9MLIrNxXj47YNwrFzC5CoGPgzDVNQ5YShi4GZ9Py4AuTcTxish9UaL0RABbTLLwKZLk
tpX4y/YRadFJH0h+4LauraEiXmBi7Dca3BHnrjWO5+yuThBJPtUlzBKlS+sU2iqowBLaVv5Q4MfM
H251ev6VbPxZ6umQWBpE66PS7No7OH8n1IsPBbuM9RljAZEEcT1PJQWuJG1Dahu46+MPOu3tG4oF
uoAjjKHWY0jV9O20aMkIgR8sppFlXRPUv1Ym3H9CGaDt9f6TnbXyZLvKgJ+uugZwrmsara0Es3t+
hQ8nItvYxWxYC5xIZSkgnb/wyyMgU9QJLu6l9xdvmNcJWY00dXKSHP7OEe4hSPHxwL5lvsoUln/W
RBHqHUngN1a1Q7WWENnplxHsemX3trkjJIXfyfiO7F4Ac9mix//2O2mMh+jKl8zwg6y7IjRq+Zss
rShTcezBgPBIncQ8aDlIsjVEK/3iGpF4izJoS0TWb+OlHN723kJwT9HepEYUrM/AbJgTBh9wB6Yl
Xj0VcaaPLg24mHcl7mdzl7CTuxNbwaAj4hD7RmGA+aKYBUiJBaQHkcw+AlAqFYXj0JYcbTdz4NmY
Z33Bw/kFyWc0is4S83WlmVzhuNWk7Y3P5+dY4b685pz5rn1mVVk8euNnOgiTG07s0Pg2pnUCD/SY
/eIzzG4s4wyuMPzxa/C/w4hU3WTj8Y/RpSPVd3WrFHrHfDwQDdEaf2+y/AAbqRoZxgKYYd1lOv5W
y71l7aUJ9bLejkoCIs9UW+j14z6xrRwLXO07ePrxfv3v6GurCu5AIvvF9Umvsp3FC2uJ0pp87Oy2
epZ7IksKdk88GMPlNuRqqfZOhlI8A3DxKOI7fJIQFDMNv04bKweYirGCbM/Ze7+tJG8IWDCa5BHl
Z7FmTYrE2E27FXr1kdoPbUYMIJnNyc8F3UhVzFveVOK2RoXnH4lLhgANADy17ebkqJ+m9/Q5/d49
nP1k+ehUCV5oqfRQqs9CELaKPluQjp0MbDWox0HSxMfjSwSc08lwyfhSnCV7nhW3QKuUdMUyQBoU
mXVGGrVHKNwkScokRiGRm4bAoQp+3eFPjLo6mxm/tlWuf/3gwsOBmUZ1dOHzu1ZQx0IILDiRKqAV
hppaD2tf2T7Wj+kUY0VMJABvPxJny0PO4njBDXkRyOOtGFNSJWQx1wteLNs7kk8EMs/zJ4U6jhEV
DCYiv/+JKJ+t62widGtI2Vel6cX4x3J0nJQPRPPkuQ7eiOmRuOIPjRuJfe9oIkIc5aMW0ay8v6Kl
35fPtdN30W7b8cdlGtceVGFIJA00W0k9sFJAvmtsx/G64tQiRYgo/5reqpu/ETrMAgHYsROV+u2w
NVMBuTRnrH4r/TM+Z/fdMVmPYVonl29fG8KK6qYdb/1UgmWorPAKVGFkUKM8ukjE25aY1FSIluMm
g6AqXD6uv0WD8mr6ILDZYvtEwcFSAJYCvwAdxb2wb24k5JhKBmqiFkRRJV0E806jIb45LZ5U954x
OaBr2zd1FXHww38WgNELGyZ+mAoAlebJoaTZu8+KHiHl6Ow9PAyMrTgBfGjLLOEy0GgSkvgAYqQO
HylAItNyoACIrCtVAyQvWtk4fNE5AOS9NqCazyimV88j56OFDq9HNCA5TpRdMOsQ9T+A3RItyah2
79Cm2uH9NlCv/2vjvrnCwTZKOSm27+L/FFKRWkyZph2aXWwqck2XXAGQxiELrAky4lSPkU35mNnV
oWXPLdNspInpYFyK5uVgvRO108TaupCt1g2k13S0hJdLykGfGjiXkLNbBfF6hAxcEWAFqmdVuAlC
ekGA2jmgtpx8kOTeQiSZymKSVgOPWIRxSiRoljN5H9xhWFzqwLR438VKAwjJpSxR4EQUWDL7NwZd
X6m2tKJv9BEv7dvl14g1nP7QHB2qChrZ/S/YkN0MoGBSbzXe7EznJfC2NfJ0Jq8b1835NYcX6oYM
2h23Q2SehKLp3CiMrhLEvBHIQClY4bS5RchI0GJKJqYaEyt5v2yvmM0Ky6v+PhaF1nuxTUg3WGp2
btUbQXG5jUSneaUhaPmotr85mLKW7fHdXABVhx3jgUG8c0ZSbz2mM6Pgk8taWWXTOkmSbkBlpq1n
3VZ1CfldQDItM/gJ++PGUbMbBczXgdD23M6hhED2qhfsKUhr1OYoKxLxLYY7PdwqSFREJZsghTdr
O4VPxGCIQj94/sLMAikRoKGnwjInm+l8A+FUJ64v9+fzygLUfYa6AxaaZ+dEoifgA1dYBuRrdzVv
010rtpZeUbk4QkL+BK9LlgrijNmWSb4sXl/SPCCwOvM3tic3xo7cUg1o5NAJ2KL//RFkrA4KQsSr
MJTYPSnY+xdxDcPiI31xNK+lhK+fMcp1BpqsYlITen61wuswNkLhSH40f0gnb/0+cBl1FueOtIas
3Bt7Pk/xIxB06FAfcCb4raMBlxtoqgjBmtyxInJqOUNoRFKfHTLcXG2qe93Tlhwyt6qFDUjrYtM+
9hJMLgx63Hx6C3J/ReD7mnBn77qLMh1PPLo+KPyVN/5K37mj8zFNlyyGlJOOBgxNiDu5BSRbLI2K
mne7xTzoFsbKfpgvf9ywGm3jwjainJQBkDfFthQXtezSspNiMR5xxT1zCbiAF1L3ipPm4kfg4pM+
NKVL2MPCry1vwTswQMevLF+SozyKxlFMMUQsgwDvzvr+dr0x1/LlzOYA7ff+PY+8ngRi0LhAD02/
Uj7LWQ5Z3ZB+8f2yIMgdPKlVSwSUyqqbg5JgHs2pd8yuQDsq+1s/edYwoaOZjbHdKlLqWfEi5JVO
ZZlc3xFlHkXdCytE6l0PpPeBMahpxwpRnP13jwqVMjGiopCsq/z14CR/FY8qXSzgU9FdKylafz5F
sBQsLbbK15tdeRDsNXo7aCSaqhGjsm5FPGJTP0led3ZMIFb1Yu6OFsK/kBJaUsJeWJ6oNoNEo3ke
hC+vz1GpvmM53Ds4YSYMrUe8jT9M3JLl+HQwPXIvolfc6nUnokL+tNBhYOc8fLQ9giGdybFtBfBo
9USaiEJac6p54G/6mbDyOBIH4qMuW2BtzUS0BTsqIRf1QhYqGcNst7DO+UBjuJAfg0wfbIOnRvXq
CzciS7vg86mMi7DG6VDX6vZ7hmdXbwAyaJQHAUtcLNRJdDoiSBTUkR9FZFq+AtLxcppxPnwXb5YN
52kRIBkeyhd5C/8/gCDeRMlZWky0sZ4gbRdaFbNoChcqqCaoCqc8/ju+SoZKXMFhBbiWb4OYLNXI
sRKqmzemqu5KOe8DUYrkAAw0ehIiLLE4ocfgfPPt6d5uUlNDuu1nc9I+4o7UY/iyxYtTl8UhlFJ/
r1LXaA3QHIqhDbytR36IabQ9O/VhLVS7tYV9zzZ2xCVHwoWMvTqdexkn9YPfN5VoW5G0gzojAjhi
uwxmrKL48OgxK/nvxQbjp52xcdYcI8gyj21XAFj5DW1IC/klUz/+U2lEoWv23xLsKAJWJANHCuam
yQr3cvBuXajkmgzSacmTWESMGEsKGa9LuQ5X1sCmtxOwrISA4PXvS3nxVLC2GAFDnsSypMl3G3hn
T40hekRzQ4OHSfYuZo0am9iWNFmun0MMtWFr7jDiMp+iIUUfgv+4Kd0oYAmP78oAoCFtASpwEs97
KNiFO1XIOB6qggK9UCs34v2tebke5VyK+hBhMb8yF6UmmwHWgpQTCRoxmSiyI6TA2cl930YV/xnZ
hsOQCGPzWQySJY0ZdiScJTgV+oUFkuJ8WpbbI0It0EaNxhPXWCw2xZTVHo8SQx7XEO/mD/eWWPTs
iwzpJlRJc0Bwl9TKVFdePf4HtjW1OFEyiPm3HDW1F7zvp+3L3RXz3Z35TOHT1/npnTy/wZikNUU8
z4zu1AWm2y/rrBIf3jwp6f8b4O+qpkdjwJmqsdNFX1A/hm9itA7lGwUrYreAvY9rmsJatApwoLS4
EYZt/VRlSlYhxDT5BxO3ZjY80iKU5rs363YMQbtgHRSPjd6wK9zCodPj09TIiMn6rr/f424hsgh2
waUUrv33NK9nSGhCsO4pzxY0Z47keyG6egFEAYW0BSTmu0Zv9wqhOwDq35qS7quk/YVl4TXBJDOP
CNSGexolfehUnDCZSal+TB6X0HBHSm4rKoOL2uEjgrqcl+NKDIpDU9xdykSRaRaPwSOHiFvu6Q7I
Q2Glgr8Bi4irq7EI6K1oo6mvyBvO07Vwcg4R1OkyOm4/z9QlExbX1XAAgYrrUuC2Vzo/unnR2bjC
9k4LgvpBRSKZGNaMpmOVYc2Ri3b/BocX8ph8MnavGpwvGyF2oeL5qLGKaiMHTY2h9yiznij010Cp
uiqHsbQt/0qskQatv/jiuOsTJLMTgaRV3zpeEnFzL1XLiNFXU6Ox+Ix0kXWV8vxxyylyGfxaHiXh
qTEl3tw/2dlFLCB/odfk/JtosQC2xvsOsV7JIUP0LTROMnWllKcNHazC2M2Ny7ZGFKTRdgdAJrvq
DF/qbrcy+HH+oeSQHj597+8+4eKrExGIyCL6mFT0ADMcSpgPm1W5hs4VUmSQE+UGJeZBzNUFHNF3
tUlyJnq283IYRXryv9Wmg+6YWIRm+v5foSFruXjoV/HeQ2vaxKDndORXN9A9ZknmOMmrvWkf2vm2
jffCH0VkLGVevgYyN49Rb+b6nKSiR0HEvDm6r3E4J3Ks/R8WdMxDrPHE0MOy1swrLzVtarmYKTL7
pGnPWAij6megc37qKcYVFaJj/zuUAMGsAgFTUy56oUwU4ZZMcCB9F69FOKgpxtQYCx+/hiJesfgH
L3Rj3erOXcE3YLsWTXyLFhOsMnLLKymtxKaI2yd17FBm+rE0/+WByar2edIeU1THnLefIb69Wu8I
ALbLSI+2YrsNbgerwq/uFU0iPawGxfeJiXYqK5c+jEzogK4WgkNfr9VPTWIdjx7ZXjX8BEBnvzVf
K61og0cuVX0NXR82Ibrt/74WABMsizIQKfSTdui3p8wsaM0VUA5LC96AW6ViYzlwDRBCYI9dlomc
0WPnpwLUGFNE3m2qJ5WS8r4fpabiR0u1cWeM1h35Ku4/dJ7z2ysW5bj8yUXgdXuL0rxKc6u9+oyH
yR8SKzmjxRaoCuE2ms2jNNHtHBO2V7ur0WQ3P+j36bHHoJExXxAQ5RWAaodRAc8mL2C5WLPnimPy
nRxfJkjY/5sxQ9rasahbiChtCjF2JzEtDfFkWOreQiEW4OSzeHLrPz++J8XalpR4xb+QWQEMpRwW
Ah9M2WJbpWQIIrtJQ/qf3IEGvdpmJuKBCazmuQQxeqYgL6N8fKLracA9YCis6j6v28iy7rC8yMuX
5XkuYQrB+GHCPyO9h3KR11LaOC36tubz97yPEp9Xo2asMS7lPvS2u39Y3S6dfHP6gzB/pDpKqtqB
hNCLX2CDUU2sPzw0NhFtv3zLkhwIqiwu9JR9kwQBNqqzuYwBWZpBJIORN5GwY8GhM8Uz/2qLf9oU
fYj5aCSegTAo8popgFNH57kz00IwYCacJXf5HYlQEVFmt+3yglrKAyy/otNkqNx7Aogd0b79mLAK
So1sKrbk5hv0UhtTC8nJhH2aSTsYBsuxTHEsgkdrA1fsVGUzjZURU7jJYcFc+W5RsTX0bhT6M1/W
yNsvXerEwhha0hWB+/gbdMp0s/feZ+/qZwPs6AN8T4abtHrG5kHukkpns/G4U9FC3h0AVLPIxrdI
9FaAXIVPywAp2KOFcTfBEM4RmlXBj7PoFhHaWFgx6mL1Y/SyGUnNlrrQ6fQRKajvtHA0tNTH0dN7
NN0CxsHd/xsYhHFTL7zmY0P56W2F+vgg3OgsbSfHeExWY7CY2U1+ZSIwEjQFFlczd+W7YUj0QP48
eJcwVmUFVGbAbdZrSWikIp2fs4471q7zcBm1OpCNzy+RLmW7kFrHXFoFiZqvVogs4ozTXeghp0/O
2Nls352YI1tAogsNFDp3pj7hBpWlNoVPWJBQZBoT9b5Z+wk5El35dfXkCT5rEO3tjkRZkPwn7760
g5D/N0mzxolk1yDR0Y6qOCHB9OTCnGUYNKeayB38MipVtr76YL3rkKqJ+/La0kyQdLIYWXolQR7l
6nLa/7RHlPWPKf6fE/km54z3HL6pZgR4zsn+Bmv9LF1WFa83vb/RJEqHsTRk1IYUoeV5yHpnGnyg
lv9Ivr8Tj4PwepdpC1rOALzUN9pZzy80TcMrTzNVkhcqCHJrevlLUmDxa3oTuANoY5rK1fFbPlN8
HE4YB8Gp1EPFCnX28UDCRuFC8R0d0zmhnp66bKgq7lxI5y1dRMsrTWeJyxZUCvUqAvmJLhMC1C8g
ogwwBVdD5vm/Dr1VGTJKMP39cgO8F/PQMWcCgmRCsDsbxGaloIxCBuY/boQmKwk+Fi9YsbpJwU5H
L0lbQqqG4p/MZEc0nVvZVJRqIDkx7hQOycXOrm71rLhco+Ggoqo81TKnLyzBV7CmEQUERLjBbekp
g5OJW95PXvDYvg5H076OVRRsaabIAuwnbdWqWv29wjVfPTN14huMEJ3SO+/lrCqDYKp8YwqMKjyG
SwctkhcvDwqOsBRDOVpmf3q+zjW0UyZ2UGVIVDCPPx6TFZnCtvCpKvoxgY3b5nHg/LeDcfpM6zM/
h6D6vYiJjIcC//hB7Ij4UXNSbDqh4ZwZ5cv4ZvTYG05yu6ocdvrWPAI13EFcfvclWuM3cRvLT+kJ
tmgS4PoXMMqAUnBNnggLcqMw7UE6TMbAaD8oXpvXvjBeX60+rie5kIic5BeBjhIJY0k2RxkIjOUt
ivBwPvmbk3nBiNyfkv6VYT2mET1JkbHhHU+HlTOOoiWU9nsv+x8541uKr+PEwbNNrN2yaikat7m9
w4IuiIKUq6uXdhdx6sSEvSfsk54jw1MFv7tAjWIhePTBi7utO4IMGoO/NadF8Xy5lzpAiAO489CH
L022i4oWw+cHX1nCOkHS0fDRnEnmqLi58EwZI7rxitY9IhAJM+ceQHdSsF6Hba4y34emWskq2Gv3
PJNZpMhgEnyhKVea4LGD+uYOQJRSXqvUDRYo8a97UIT+IYikq7xnTL1vBqMmP6Clp53II5H187Xc
/xwtxZDc0gP9NMKPXDlamNyanou/tk49JwrBXXxz6FE3sbNdqdw85fXagvswuBLcN8XgjNdOihs5
yCVmRzTAMtMvVfWRiReIwKXVF3w3IcyFt4aUHinRq8395K+zwbe0xtgopLIP9Nm9qwVkI1TarQLV
S+OEuiSXdwkXJKMBm9bWNnbF/QsT3BlvhHlogSfQgesaloUzfa3DvfU3QdMUkwPNvYZq62GNS0VD
5sTmY1j/MI9ST6RPchkY66A8j7n9uHG+5NbVKSF2SaLgehnLV2GUoLfN4+vS0sZXUsgKNQndpBX+
7OtxGDgPUbxznfwrOruZlbyYrcAdHnDJmfQwu0J33hGxdBviI/kOSSARu+QD/co8nnB4C8swvcKu
HKO01DAEKLlVkOSiTvanGRD1GMgklPJj7aBUkdaZ8Gs01fIOALcl0soVfjRLcZMhT8bA4kPvGSR7
efpqRs5tWFGjzdCfh8MjjZO/kOC6weq7EzAnVC71wvq8RPTWvDh1Iprxusxe+7nctjtCmgnsRCWt
/0wkKQccCwnwsPzlG3f/nnZfPSbuetF4Aj17sH06Wl/r7dcJV5KbIAUocd57tOU0F99sK8tIxs3T
OXbgHyWFDDDy1sUKpm0qTgwQn4fiUWTf/B7O/oG7DSc7wJjoMhQcQp9Ba1XnYflQf/K/6gjZKlg7
coRGi2yMZdjl5TTH0nisILFMoXA8ThAh2s0SO6s4OyiGLLxEkwPN2v1ySwnHFc4IXj5tFux3mVdd
XJ2IIEfBm3xBxYZhXPQcPIiaLvM7ExkHQVkjZbgL6JqDZ1+jmnP8DObX8/hjJN8ZU3X4vvS2lks5
BuacTPFfL4QBnYf06W9q+AGb/1aP2Z/xJRFOhmwAbQVT+OUsZhUl4LWmZ0CKAaAKD05ggKog3FY0
Mn3zE/TWuxktzDcU8AOaMVKjnO7D0jq/R0+KMqFqoSZ35oCCorVyqT7LLyX2hbY6HihmEkpH7507
LEyZl+ZG6f4LAEm0rtikpiBDvTzE3CEYy5MMaJBNdlfJoBUaeZbvMV4W6nnISh9IjQlkMNKKLPLl
woQ50hvImU83wO2IYaYnjbnG4DdiVm+mqKwYf8mk7kpln5S99e6txnUArDKLMn4e4r6hKn0Ito49
VaHhSDnkUel8AiJOlQMnSTp48Dh4g7IUk6UxbjCgoQygPCTtfmYyCzN24Rhjv+3gMXEc3kpfGczo
UT3U59aDrPeN2vN4092XxTPiB27xBZoXoD+qwi1sNoyYvXXcjP/IQUY9ITMZ4eVaMEMvfKw8SUIr
tDo+wQPRAtijFHQQNI10hwfo5RsQGOvnOTqIvQ4AZLIsP4p4j/ukQ7QKprnj10vpXmv5EO6qSzKX
Ww5DoJYrMMD1IyqTHf2ZXshoorUas8QCppzv9XG5OzKkIXWbFTc110Khwrmd3KPi9JgDZNpOj9UG
Nkc+zbh18Fc+/go2IHJL6jmzgLmEu1r1tkirVDQLjfxiU8Jtj1KAoXUUt2UddRxH1MvxHijBU4Yi
ToMvVpG5XBE5emZbZSgSb2w7rpgg77f2WRYD3kRtAvybeodJRCXLCQYAHnD897daPihFpIK12Qzm
iQJ85jOlA8unWynQ8QQ35ADur9lxLGye5s1Jy0UL7aHZcwLnnlRooY8+qtqq9E9mgdeUpDBChjuN
f5GFd1q8cN+wZUoDMp5qdyKlmr6gXXE5F0qYdABiAF5Wz6BqPQtX062VBleXk4Wws0zCrpGstEgj
ot93oF/QnVxdnhVuqM0yfPKXwP+2dcQaXrp7KeujHmYr81MlwZk2ZDBOC5UUS2bwN1QHBKIN67R/
fl57E+/ZSbHfLJD0IPao75UToHOOY+gWZZUH04EDOFnxx2L/DcUbESOUmifmLB07toRh6oB4VH1P
4LC3VXkQiNtx7LBCmXKx+mr0h7RHVUB/DtNxo3euwjucn5/Z3v2MIyoQdMnp3bzqJ64ySM64MBtS
Vc/xn+fCT7FqVQAfzhOQ5C6zeR+fJzIN3RHeCKqBXkaKNBsWwmjBvIfqPqU6tQhZN8F/zkBOjw4o
ajiVwQVPBCv6o7ltGHWM7b9y8nlt/Ii7uslMuc/13Op9tMbb82GosLpDs8FmS7GQZOwkRQKdSc1u
5ekYWBpSQK/qZJA+HuR5N96sm3P+x+uF9XB0x4to+DIwno33LWLDKVxq6uJqXOb1EsxqY/VdgEC+
9UMW9j5UjhlKWGuSEd4mD99foI0W1/BhEJ5rWO6dNIL8xULi2KFBwZSmyVsel1FeXzajkDA1iNHw
zwURn236QvIbRn2Q8pfD14sWogZ1ftWugT5rPN6g55dAZmTp7qFIl2Rb3vcESBbGZdIz3Us/+9zj
pH0tMZpWOPH6ER2rMquElMA8m+Rwc6WZ/GDACr2gWPNWBHivR1UA0MmIwYp3cQQI/Z7mpaSLkUPN
IKPTS/ev2UEN/Bvn63gj3aWidDZAqhoL8c1XwaCdDcQAfmP9HwtZvz0OFW82szD8AeSL7oRRdlGE
d7HFSi17AuZ1SqOEwfAbMAqzX8N/wdUP29APqzNrLzSzy9+w6jexZhDbFOvHldz8xSIu8kQa+sjO
GPnGLruUUM77FfTicCTnMsFGIQTzWIPw/m7gWDXObb40wkple+Qoe1Il2PSc8XolPwknp9yKBtRh
8377WMvaqmvy9pY/CI4CtIq4M22s8Vb3SwtXpzekZeEegfAx7P0S5ZWmBeVmc5HGCkyaUz7Hf1Lo
2qcvcOkd0dY4wQw/VGxWPBgZHSgtPvPeC6buDUmgqWstZuRvaSK3Enrbi6Dxp3zpvuh8gNkS8rZO
Bhl+lhXpra3c55ue3UGPt5AoxDrl7SpGSPEPT26yyvsSBgGB1PUb/5JvL7FtUJ00YBDjSoJN3Meu
GMYWm5lVunGFlZu3iuhIjUxop24/Ki2I0duNT4QjASEFpHCHczFReLItt5YxPABt5DzVsgfBy6T+
zTVbJEsblxfMq6PC/oVv93rCGtoW7wd5f4WuTt26k3HC9/jW0cbNtHpUTLVHieJfhMiqoctoTqIU
HyH0FwCkMxlUXeEX9EkS+vO5d+/IWHrtVlv1kS34YQOk++vmtYACU9Lcx6WjmGbdYt/YfvPBSkZU
9TwDI2FZqkrLGlLh+EuzqbanxxxplGV6vwyeoZiswRA6Pjs+AUEdxylQmHciDn+dYp4yrj5Qbfdx
9re6dol30f9dR9APe3bAagp5wyBeqUZWWL7WLeCfawXvlHc3IZBr7U0+qKZ1tWoTVerszoPAkyfD
coy1fLfVQHnggGnR95ibSwVhOu7w0pDQ9CQTr4C06ft1jwh9uxhpqrOisbMNgSLGl8koGvt+c+Qv
F8pcYZowHFuefOtY6e5taUubZbVnsRjCMEAFBWDW3tLVSRwpTkiXYrv+Se5uGyABJXilIAhusbIG
Hqkhm7REKLiKTrQwMZUPP7SeKvBqPMp+u2hVmZ6p4Nq4PSFWxvt6pxjuqNPKFPr90HGgmKaGe120
a1DTRAYiESquTjHkI1ke/xkkJa3qqUEsFU780riq872w8deVDOfNeDdsQwW8tie7YAIEQ9sZT0dq
/5q8QcTOGIidR5AK1pVl8tQYYnER2c5V8gM1UV57cDIErbkUFUF/SqGmhFIiTYjTgjQmnLg2QgYR
ay+V/EL6Yu2rEYFW7xdK/8BcLhxZbaYkfbxxMDlTM4KNK3V489f3DMwcOnhhJTufBkpJXtq8+4E+
EBwYt6NS0IjkrEDEznjA8mpqFfclywdd+kFkkltEbtdNmCgcp6k4A0QBUsBWKbIAYlCxf00cu64B
/8L4Qqt4vBdhBCNYGuTBeSrY3FCaJqEfk9d5i360kkgGMpcg1Q4Auii2M9f7YEynes/WA6iHxuRL
+hUfeT9W7EC7RnTd0hDYHdoQGlVz9292yt0/D8QEsa1V5H596JZ+RnsMj5K71P+1ewQRvOxTnPrV
f2EZaHVJ4cH0uuacTq9ZDGgYbYhIbRSZhnQEyBrzosH2f3b58wE1tSHgllruMCq3PQky5rrL7er7
p/XEwWqhKEwRyCGNNFchZYV/bJcq4+38I/TjGAm0Sbzg/WM8m+VEwBlEbeqqLo3P9Cv0vOltUfPw
uFM7jYwspUWv9LsNCQaQErdh6aw79hFXFkllK872pSra4e+FvDddGWWETfKdXFQ6jUwu9TXgjvcg
V4/k34BqIXbHEqHlW5+7P3DiRtxFrOK9tYYlX+MTEdXOqwNJp4VSSpCCA2OEMbr0t7kcRFoxA/d7
fExI7hOYfHN+UYGgejphw7xPwetbPIBzOQ47oOrRezd+rWDINwbN+pUFjPtwDljDQQxoN4Zwju2Z
N4+xsi82oEKngEn+3c0Y601AaBVaPW785lZ9hFhdsxwtwpkeyYDTQ+fD+7JJOOSfc2lO4IMQIxVF
BUKCHrtUBMSh2i/XrDXtHs41wllvAyE7wxkQNRTs7V3G2pGDGVVJqVv9WtZZvJ/Pp/x71xTkVtgA
2kCUzCnbGe05vHZsu8sG3DUcQenxykZ1G5y5SPM+rza1O6ZcoFCgBOpZNapUbZMfNJiiTwqXRps1
XRhnhyDO38zFMeQaVrOAQIIXvvRPMAb7aM6m5BB+y5FV5QsgzRp7vy6o3NFQhRJC6EtTP5CGGjas
3mlqTpIlQM0ld3yHD5jD4Jei5SM6VqrTvd5gmE9pXTEB702ApZWHYwuQ3XtPozmfn571ggtBrr75
ViNUfAkVKQPcWWb3UxtDTyz45K2eH3+ItDUWuxKiBs3jMVocy2nptOPaKCQjeunu+gUNPqI6QJwJ
l+u/BTokS/o2/IFdXLcEbrW5WVHbfEsKdSZRgrwL7kflDiNTKNsdYwIPEMWvsE/bTuZ+b01fpjE0
X85te//NH7Z2EOf9AjmJV1Y/2anVFy4c/jS1068ZHM7Dq/SJsiNdgtTX+Gd21ynXrUqODeBDdUw+
smvXWrzjEa6/1mmq9gXO8hUFRnwkDXAQobW7JoUXzl3FzMCUIgVXstUU/JOYkiaPGUhjKrzw4Bq7
rOE8o7pAQY97Pa5/eNHRmpNqvYQ833rzd9Le6qY0Zl6oMvTgqxwqRXuucohBuyKEPrjzCD9qT1Nq
2x2OuBTL14EYEyiJUenu9mnQxDzilqaj84s1WteCH4AB5LpWvIcuYXGvDG7W7lZSB81E0oNNsThr
A1MUKaQI/4hVRMn0+yp2czazxCCLRw1TpfJERNlKzY2FqKyPBuhqKHhpSn2+VuHxx0U6ATmHGD0u
UvHrSoEcTEo+0ElWayexE+GeAK31jkFt2DOhcTVaGFdmmNbe+lZC09YBZsu/BkYJx46YsnBKQZBz
gta5bC1xZ647j/t4virsuDlRi0KZVs9HX7c18Qj83fCcCf1qWs7ZuC8Oh+DaHjxnOF6Sm5W7IidD
5gEehsO3sbZUWO6BGDNLMUmYIimDelB/8/pJ+Ex3UxlOD45ZJxrT/8AzbcB+Z7YS5cH2Y410eJ/4
J1WH26zqdOhR3hHFHd/9DYd7CpGKek4vaoodFYkTqRe7WHcFkvUsiJ4KT4cS4pjni6EERhrhybKU
gNWPkA+LGKHDE3kAkGszjamASEmMbkwhpczYBOY4oP97rOTpXUKZVphQbv3aNbzHzEgsB76RcEJh
p6n2X++8EqDVVKe9VSSPiM8P6k0i9w4FS4ihh/IsNMZQVVEoDTsYVlFpIyBaN0huOJXeInDJzCvG
vNyZENYEQi/JuOeDP3k+DgkayIaRBchb4+hH16NP4lmLLS5c3cAcEu/pDarb17ArwA2RocJrwlxY
03EhcpR9HGclTVOkxcUKmxDWkRgoowUgqx8c0U5LED24EXsMMSruhOiyVBiuYl1GJTCFXpN/OBl+
oZ5kneM+3gWNvbJFVY7g1Tf42CK80kNqAKS5DMloNP9OoCE0dIomIoVQgO2TAR96BguvYYwdyOA3
j7gfYFxTO+tYpVKUWm1h3F6JVHukNHv91kO/JRep9Fih/P4XKMSg9GgjqVvBI7XtR2Au0skZNsDT
bmPG/xSIqirZDYXjB6d+6HY7MbEFS+9Xxk+lK48Br4opNBXJdAIVudMps51zRlwpM8k+J+4jlgWK
Jo9cNc9Q0gLzsYx+56C1TU3SBxv2KIPXH0uAVnrQcRIDX1y7nGOh19kwHNLsxxr6DKYRv/kkV5C/
vi5yuVRJAjTXa9a+NNuqCIyV237x1ByaoiNNASbQdee9DpKaHQnbwNjDlrrBNNq8e5XSn5BBCYrt
92vzjapTlZnhAdzaDSpEX+EAtQrkZKuYOW4Ljk6I9D3PCUcj4dfKv3Xe5Wbf4o/rfjHCBEhjT/mr
Qp/pAl+cKiay4du/4c4xbFeD188TPb2X/Ql1CTV0HJ6rTEAjsIClyO/sX4VYoeBmoQPM5QNMsqqW
0TRlPJ7z1Z8NBBsAk3tnvJ4HBjj1ODsqTAYGsxs6ExYxoM1z3QUmoVXvSltceMtGwNoWRAT32PO2
0UEXlWUb/AchBeBG06xE8DOzqvG1k1EYNbb881KrNLIyHyxFXU3LXsJrD479BtvVCH5SFZxU42dg
GSqpqw7gzoRKPg3FajRJuAI/yPgWKQstJIhfbr5JxTzJ68nrfGHm1/feQgodtlDI+vZZFVsPeBMc
pdVDiFQoLylcmBibDPT+bg5FEBqtmWdiTbm+OmDaPTdtbXtx2K6Guog5iQKgirN/hOl6eyjo7jBj
v9nYaroHEw0MJ/5jDbe0FBcCLDTx6N+/OPYywuglqc7zBYla1FmvzL5czNtHp8pPQmJeaoDigiTs
qWd7Q3t3ry5lvXaZwNYomffn0ZibMMxXDUlmq/v91WWKbZgj47MocMvcJxftujXU1MKoCAiArTkz
85qqm2dmgS9TYh4yccmgcZ9X43huX+M9PzvFndINTfz4qkFu4/+VUVudSUaN7LGnJK9ImFRDWCVi
zxOFYNCBJoHlpBoAxOwlm0hdKn4n854H+ZxYZrXDMsjEdJJAwLe15QnF8zkjxpE3N4jfLU3rq3z6
+zAPk4nqkeYyWBLJ9XqDSfqTzAjnaQgOPrSAfWPCd0GgPbL0mJVoXsBgxGxeRQl/fNe9VuWlSf70
QBSvtuttcH+wYVdhYtduWO+294dPLVZ48evjp6Rxg6gUJ4iCbE6fuLzjbUEV+XzTcUxeB1da+Vvp
8xMqfijd3i80idFJ47uPoY5OtiYNf9VR6XH6fNl7jmMOqD153rQfgbq4mH2WB/f6GuBUxKPArcnm
4xK0PLRNTz7wLIl4ubzxnNnSLMLIGcKRvYc6Ji/GaUBleFeGfNFqeiKGbIV8ou0q64Arlu+h3KMh
ywackGIeO+OrLka7WhrGZFQyU6qGa71DZbe4otSKgjcj6IsrtTYdQKpA4SvfVAr4SEE7SgyKmjlw
lbsf0wYBkW6J5QjxoSWJ3rPyUQ1uO5sR6DJ7BifocpiGoGQFUTNFlnb4ykFTk2OgZp5q1t4E65iJ
ocm+CN4nKCk9tlKV6y8XnSUTQz7yxpXYpVrkctdvHgKtdC2CWz36m9XaA5dDOjTpdA3CkHcb6QxS
PCmcwrIvonUH827UBrdGO9WJT0TfoEK8XrDlR8C7aw34LVEfXdly8pie4IPDUcMQbahldUD4c7fG
Ks6Nkr9OMQ57kbL7d6IXRwIkCMkG0tFbXHPeEr60Gext2mzblciPD5n8aPb3K4nvhucuyHmiRD+s
U23SOTKRGuALBOc9IfNL5kdI40IYARhZrNJ1b5GNXFteB9HnCEQIzhl0Xks4v+smpRaySfNrgg7q
eaRibYI/yWTin+oBuz2DMeLFhiR7k70jrp3pJSvmXEY2mtVL0WaFPVFfSNNQ34iJ9fGUgYvDhZ7N
DIsOnAPdbMrWd/f6ZNBVBgoeboL9LmySsu4H14JND56EEz805dGy4XWZVhWZofNpm9eClqSf5Zdt
HzsKEXL542/3nDcnukBujMmfs49aVVz9gGbdW2P7tHql0VPHOnqwfswHNl80/0T4kgRE6KqHbfIx
LzdOb9PtNSQACmfhUGrAGGaOG8RHHk+D4POuClx83RyuNMKXTr2JZXaI27LHDcBh1kXUrr90zNOI
JdEAW0jyIl2pdycrCxK+EO7BI02cs9wYSge6vSiTe5Q2rxSLFIBTkTmFLpTj3CYrf+MXPJ7cRfg+
2zMJ9DnmXliXzAKaiHPV/0a1P0EUg4UhR8NIxUftqGO4lFUKiHbxOHNemobg8IEn25cSDxJ4qvQU
Q6fElaIIRwrwx622/+PL+n7e/bFErmYksywOCfgNE2IL7196ms2pE1EZMYqAg0HF+CwvMqwTpi/R
i3iCl6p08gzeeEUdhalnHZBxMca9eabJVgwXVD9IZXvGe1zMFtoll20y+5qZFX3uSzReA61ylrzV
sG83paSLTr1vUl6ts8qtpN0Zp2dwA0xtu6PFwJezcoESNV/u+zkEd5tz9uoeU+FjZJSIm/SdXoo4
ABvgHO0R3HqemF9plCinVST21m4UtXWY12Kep21emQqzH8WF1aCrJKXVG+iXs32K/R4szZzXwCBR
5KLLRJbHTRp28i3mfUfF6xRw3XyDpU9pK/iyaGAhTXWlUJYwZqswltj2+j9k2ys6dumTQKJ5REEk
75DWvS5VTTS26x62BW6Apm8nzNYuBcxzIwiRRDGgf5ZXhC+xmJcipgpIcIyvxt0EbTy7VOwZOiEz
tmiSv42BoSQIW1eL1Q1V9Ag6xmi1DrRkbZhkTnIt65t7H2WpSfWrasiKwQIU4gCdKUqujvE50dEW
E1rKm8H0vEsFxYorfGw0mmGIl4G1ubPkizmX50OLeYi3CFUJ7fWDnIYGOf+PtpqTCKoFxWxlXOZb
88HTwEMCi6+p/WGDnhixOztBOwjIKBfh2w6DRILfM8iLXq/K8JkKgHOOqIqARPabJ2jEkX7XDqk/
8LUJhtvDksUk+e3+Kl3b9iA8TPDrfTuK9xkZLnJ2nRFYtkkpm0XKnJadTfv+JnbVC5flgjEoeXTC
XoKNFMty0mQv2E3SaOMr/r37duRu4LrNKGi0RtvdkX/7S4V2b6oiGdge59TdivTN2vtbGjRyj8Yi
gM0nG3Qb8Tn6Zcu6Z09xkm9t4OtGEO/54CHNdFPTiFfvBN+z7waafEnYgj5A9mscRnVjCAjsRqtq
WdXYbKNcNOMs0aRmgkYUPaA+s2CiK1WBV1vXP4FQ/zVwxTvaHyUAodI8c9hv/Ths3ALLIX/+hDK1
IfzwcCtbCWXSNmiaUm0SyVqj7x1F5l9/yzTE6cagFm6JnfarmZ9br6aWzmaByboe6QRS1Sdnxf+z
h3+5Vsnc0DLxXU/wpWcCoxRzf0e7xaV04oOtLwRSPSIPiOSHqJONM+MDsPWx5s9p+Hh9r7788SUI
dJiRmwZ/ZR7Dz/crvLUCifNPkEXNXr2Nz5ZCTVDG4G4tmN+6vbw5srhqXye1yektgc2IRat4Jdkz
wsTVDPJT4JM40Z7Ut7cxXgjhrf+4C1EouiHw43+QOn/gR8Ou4m8DGjXE7QkJpyWVjedL9BNihuXt
fKmEZJCB+7K67OrjyUI0yizzfkIXNJIzd8AXRZVu7xw6yZJaXBrT1U/Say7M/gDDq973Sg79uusi
+JqW1/FCsaInGotlSnxJ5XYckPuRIn6viY/lRGZv/Nw4VR2fuqW3BrgCMN0qmRNZYu//418y/qD8
sG5IEKxCFQbfSP6NQ+ZzanpOkqoVCxvd72TWFFyTdjpTxC/uYR94gQnYPyq2+sFwtLipF/3e5VMI
9atuj/78ykBgKiWHfYm7NJSIydFkJr9k6hi2fNNDtOttThJ53104FqnG5BMhu86laa9ZK0PtmLRW
omLsftJu9S4vm9bsjXb2/YxC+ijIs0X3tscUBfyA1R6V7WqIorOXVGbhJOm5My/VYGPfZEZ/sQBl
9mL/3Ht0arvjqj5eXwc/0tE2ViWjNu8QqNjZbbRCBuswyzbnv06hpeQysKCuQcYGD7CHGq+kWX4n
24wnhW8e/hZwiAF2cxGFzXHoRtdKO08Igim18SarRfeCZRp+ov3QWKYHiqjZ5/ZuO4M3m+8kVMSj
Gxkan8K7HrkgPlMHoTfSLMa4W3DJDg2bSMnoMQUa12mzpDfzpBXuSxZQAEqOrnB70ZvXd7muJI7W
VkyuqBSFMsAlF0aApi3Adz3DUnZqxudOktkKEZXBd1hLsRGch7Ty+V+8AXVVtSVlKMLpjFudw7dG
eu+XTcxqzk3n4NglrF5pC/iAyRq+BMHmdXcQ2+IhR2JjW1F9DrNw1WJXjX/4jkIkTCB31BfuggiC
nPTWwGmeO3lUxBFRZtk6Vbk4G6zkZiASYxdyUxtnTb350mIffBVyGzGAIFLvxYv4oXWDwR8F6AA4
XqvRwHdsqvoqVa6bwqzcAh4J1ACvJTQhrTCsSsZJZVuWLZzkytoKvOn2rvF+eJxqUYOF/+zV45DF
KIm/ZMEovWf0wKYrarpIuNmVGVRGxrOAEzZLGA5jI4GeL2iwu7fDlXz9JdxTN3gqgOIN9biYbRw+
69Fp2eG+pR6qxqb5tIDU8G7goJ0Uey1uuQ5V6DkJEkPshPSsBYswfQ/wmwMyRZlHZn6qGX4D6j+a
e8HSirfTNhfosF4E1R68e8Xj/dYxw3WcdR6n/TY5Vk+kxNGQJAhi2WHI3kavVL6z+eTyj3Gjm+RG
Pz1f0qNxbVpokqL5yB9MlxOUS27Pt0iX2/KDgcnoGfl8YB5GVzUqvo6bvdAlwSFKqFstsrWSqYTP
5mnNXoJsEzwPKRBTvEwFPuK2bJMpfSDvIjN4b3LPJ/IDf4zwE6M4jFjmWKTbc7Yd2wkv5DNvNDJs
+Nqzg6igVe+D3UQQo8nqUfW5T7cGUO5C5JjXmcyeN+l/1Bbq5KsIFcEmmp11ILurEasBF6qur/r+
3FX65oo7qhj74GtTpEf4NMGfesHjcGDjH/BbEQYtGj3VvAJ2haAxl3c6fa8tPnmZhjKhgIcAQ0My
BD0HwtHc50WE9l6SpyyiTRsm24e37UAlykuE30WX6Lg7myWxbmqoSEA8Rqqkh1kk9CybAHl63j1F
d5j7uUhpIbl1RTcRZviJoZX9v+zeXmiw8FfITckM9c3cOrXtzMe75QJotxGQJEEH6rCKiUiufUB/
elnPrpn//VCKw/dvmrq9tHCExCkcaAG0paxIKykBEJ8JxpJySm+5z6Pg/8eyDd7qWqY5fUDUpBEF
76yq187ZeWEWx/2QBbEKyB1h7dBOvq36G6+3hBRglwgkQAlpvStUix/oYQ+e5LJWqEwPRKZKswpK
5Dp8fpobVjMYB/n0TgBF9Yx7WkQodg2Dpc+eyuQ/dicCGC8RlRdWLcyAKmdo7D2aXUnZ8Q30aYyQ
4FXPZTA8ui2/atA8uL7xRAsptg8YQOwMUTaRun2VMVREtjycYZhX5EezlV8Go9DYlIVY6h47ofEq
Fm8qk2mQdGyY9c3OuACE+hEqWmVdjKDLWO29Mw6sqlTFDJjM37lFzwonPvCo0jig4c8Skel9qqun
+4sfPKppkBuggj2en/H8FT2TuuwMJsgFQWc/dmYKYQhC2Rode8oCxCdIxhZgU1vfTILE0rPvJ3TN
mWb67mHQsJ5IlGot25dLv98PURBd/AXhRHDQRWHA8XfUkyRwKO0Iw44v8B/wVqIyX3JJ2E28XxSj
lZG68brbOzRgBImfwN25c8jhBZLbiVtJdwpcos/k0ptVbEDG1+0mjZxBf7Uz2e/9V1dLa1svh2JJ
L+QfW02D/XGpUBE7CricC52YZMWnWS9oA3sczX1IUQ0j3nc49NwGjgHiX/utnoGCvL7Sh2RD+HtN
A5eTZmtlMpAp9GLT9lz0NHJbEzB17HxIeVgD+KJ97rPl8eatlbN4H5gzpjpuxd6BcukZZ8tCdJgA
GVpq2BER7ge8dTo6tbHl5Ht5m85GKWKKT9RcCdpa/HiFzOpWHxWMp6EhgCNjDy1T7eXq7cPrt2m3
Z3YY0Zync8MJBa5B8VFlBa/aDucFkipPZTB2hLc2JTLeVdKGw1kfdHUZ19zhCy3+9tCSB42MTjT0
7G3Z3ALeWYMy7BziPUf40TiTmJIVxeUkILfhJAX8hrKILGR0gbIm1PRjMDTv80skjPCIjQaoIdMo
KLfr16w1egzfWg3ty69Un1qbzbr13wNTOQP2GEIMaHxSqCOUY0FwDj7mwCvwk3MLvmkF/BgpQX/T
wblQRAqgGbx1ONEKLVU3qcALjqIExRXJ5fYaoP1qrqR/VdUTxmAqR0Y5Z5xYrdsGUpLxO4vD5F3P
XxydprMC/JWdI4+8SWEzL6MSFCT0dl4a4LI3Vt2EIob4qyiKwuGlYUdDqRKxziQr1il4Tg7p5ydf
GeyScTX56ADz0oYzld2nx8Rb+BqrZBtfEWZmMtEAbofidog2YaYQkXOR+ayZrU1mqwwGp+grOgZi
8KvnF5JLk3eRv007Pm2Y8AUXs/f8IogkUAwCBowfKkLEr4EacWda5C+o5GuU83yCyBc472UACqm1
JtsI96JM/tzdm/lMAv1686AXe0stl2NTvEG3sBpGb5nMfupZdCewQW/xpe5c663vbj3g5+TNpYsX
1KC7XCRLuxotjpzZ9DWpBnpVPJX/1egOIDjZNIOfxGpzBTPw2vwJYugmZOJNDQXL9MNo1zlIUV2Q
Rdsy7UQwe7mLQyDmRjSGbBT33rO/rUQHS40lwOMWXo9dSbQLptzSwtT/oppJ4j/FjB1wwmtGnmYj
DcHb1y6VR6Z7+gZ6yBORmGzlhZEgsoNPLFhO8s+bbbc7Ms2oRq+NXUFII48pj0riBSMt77GGuMxh
VnTLwcE39Pt/4h88wmoyitXtqLfB+dVJYXqqwwYtlVW/Og2JrqVhWtNAXTuPKX5JY9dUWrpfUUPj
P2Amaqm8JGGYK+71FdNwmO00xfiMOTA6JD2tYPE4TIRxwckQgN6ZQ/cIb736GCKeg/WaKwdXiLva
G+RmAuCmoFNjgENu86l00AszKbi4fhAhU3KSwMVz571jarskkbY85dv41Bf257nGB3FYEL++YOvi
81SdVFvOegAezN4HukwM+7ULrywKsT5YYzCbqSjSWJHO2sV1wrz8QW28cxdl8oh5wRCor70Qo23o
SQ+uVUI0W2HQqCl4M1km86OtXNwD7byC4UUhdd0EDQcdTdg3ArFKVv51ilFlnDgsz/dSMOv8/qLD
8+gjJnkvJaoItpZ2mNnf0XUcMgGrrf7UecF9yMdzfxEQv6taLmhnkkh10uJ5V3Fh9a+7uHSRV9Lv
3UGd2/D3lfDWq33GGHCXmMnT2Aa0+lz4YuYZhJqOBZIQSPDZZD0x9FVOdC3RF71DnB7JIkm24P4V
/lJRNvu2zdEqwQ3W/8ZuLC2IOvJNoKYw9p3Tix7gZYCamzIraRRy777886fMdDn1G+JnB1JU4Z03
dRJxzflMs7UBa086S96xmEQT3OlRpwAc4uipgbzMlgPY0CZ8+/w3MO5KO6rPCqOYlvNjPWBf4+4A
NOLTRZx0kjhszfbl7JIHWzlLsD8icEly2e6PNnu6wNoPz5INz25E/yv0A6mgA/op2dg+oDNt2U+S
FX8tkB5EaDZsQgtDqzBAp1wHD3lEpYvDeWTx2Yhkklv/cTWhmG06UlDHNqCxy3nm4u5s17N27555
uNegKTfQ02jAKUK8Eq6g5faYUpnDKJyZubj83EEUltf8agYDb90x7LZJwmLgjJIekV4eSACbtT/e
Oa/C+pNfqF4X+e7iukBDhKc0pXkITvUHV3fl15tWSU3eXJwSmR5i2b/1fnFaUY3vFDibSZ3LqUfj
hE9p7uRxY9iPsIvIv4uX87VRzeJOlH6si2LauNieR+Y8x++5vFyLGMdQU5VFE6PWF4aoi12v2Oe/
jeBJM3HwgJlZZNp229l4nGQpPMlPpOiEFJDGaXQZPDsEOJVI3X+PBAqFcblq6hND4rqjNVao93Yl
OaW76BPJ1GEDYkFdrpxh4wzn2BLAN+Hm2gO1PnBQHTKQjYCqdEvBVoDo7DOoYTe2JWB+5Kdev32o
mDJCBYMEazmC417ko8UC6Utvm1InX3OdEOJFzrcY5iA9Vwqw3ZVoOm6heOt0bsQs+fj24RLSC0U9
50t6J2xqVUQ4bGU8/5rn2aLzAarFHeP+46vKvMfsPBrMKH6AU20cCVUqNM40Ve6mKkMCm3olw/wJ
FH2VxIzEGfv5EGmp8nHfXWcxyq/dLZYU/CmT6PbYWz6NkQZlIctlSm/ZQOaubQDqYr5vlALZBea/
auIx7aW7xt59QvP1coAJ7GQ6inXIFuQXSLAIn/1PN3L8qTWmcLS7f4Fm2gN9LPbS3t6s4G94car0
4TZEX5PkGOsc0cXryVqqMogxHHttUoPefcdeu3jWQ4CpC6v1254ANCbc74wMA2SCsZ6SdJnbMXfH
vJZ1BKo28wE5gCqHwIM2YglF2AwO/+pbDcOfiRAy62Q5Llaq3jizqi+N2CTqN38qUQtql3D3VnlU
cTzK0UUO5xjToQmwgVYDlUtOAYXAk2GZh2hitSKCNaseYj4bZmL8BYRqBhrBxM0aQ+E81TvstDTh
caHbeU3/gB/41mFcZ++FVQ5NIDxOPLpaAaYFV3zzopG/SvHWfP1b1FoD7RC0aXuA2pEcAk+x7f85
OPrR/cIR/wmyrp/M8kdXe7UlsPHKIDOXyAJVCWaC4tUsWH7TnIrsAoVfzcWnX+J8jYalkd0MeetQ
pIg4gczFPhEWv8OZRPbBe3qLdB2sdAtCtpk4S8/K2nuw3jYI3BckHI1RLv74UMYljmDpwyyE3uEF
ygKN/zuLXXCQmIGn7pKAtiw7oWwhdCQzUnquAJibY6WzKcBw6XEv7hu+jbcDNBh4o/whTua5ZG8Z
0OWHuov5P4ME9/VCli0BPsh52OaNYbFOzIrw7JSLZcJ9VNCD0XKIPMh2KnWu/sfXUmK3UUgJtL4C
WhschJErRZo+wH2+zL5a3nJk4VEC4YyJV0ezETiftX2ulTCOiPPQG9M81iH1O4Tek0UCCu+9Q5P2
Vd/77qUkZBGfvXsIbqOOgdbQ6fM28oxhlmnnS2uQt1E2oD9DD6viYORL6W4s0SFqEO7aPbCF4xaS
I7AzYTi21tUG5HHq4N1gDrhJQnhDg9zXIa42kMFv/pE8uEZMkhotJW9F7/0QGSIipKga6QSKoWA6
uEt7HslleBl/0zBRbGTRsX3077pWBzLp4FSY5gSwkTJVNewuBV/BtNIJ3yjrmDzGXki5p2mbZe9m
L14jTMmTQZXA8iOhFbSIIaPjiYHNBX1+OaxKtUhXej2Om5ieMYg4XWDiXfWFG6K+Pw7zN9Bog/bM
VERywQoW+GRXvJ60zywXlYgnV8jc/bynO6y+mZbrHe0rEtGtCT4pNkN99+b5yHbtczjcd/NbINsT
TR3u1Xg6yCmsbYlniGNQkt2VUEBt1m5UEX/Tp7s96ORcKu7RVpCsoJKLhyEpVMwYvgQOAduT8OkJ
zHNRo6COhfReyTF3s1WzEsP53hTYTx7U04q2FJKelAR4JMh23NFe+ZI8XXnIkpUJ48NCsMKxtQ++
CLY03Z3c3R0+zqesG4CvjavRNHhiBwlH88wn47D1qeyaoDApd/9XiiWwJ2gAbX/Y98B892tjxnQR
3z6OGYVwtLB7eEBt16mS2WY26lsuci+TckGZWjH7urrHNcySdO1I03zUImcdvKf8aWvAnwkjQSY+
o7ZqX6T0qQdeskNtqyBmtw0KBndnrT9Bb1rA7H76lb6iutnzgVmb/rqJh/7Eey5YMHRoggaCt5U1
AdKqBbhD52YTSxeKiCavSlnqy3JyQZ5WuzZhRSaUfHy8THVTQ0JGlgSjC7p1Ohzv0VHLyc81Ahw3
QFlxAxVgAfXaBuB0lXmws7cc5Kdam7zVxgi2JdcC5ZWNVJ+4NH20SkE57uB8BJMZondWGB9sSWl/
KiIT4mzw0wwgaynrhpB7+b+AlZQ/IciPmV26Qs5CL7BkdFT7gY2UTZDilhu/O6ZCLe3UmTnWJOES
m/uhh+NmmpQc9buQjZT4a6xl3kkHiuCCcuyX3L0dpiJCZmq01MAcKFNdxa1BNdBrjfyTb0jFPJ5b
XRBfCVkxiiX8z1YPalYh3cwnxUREODn4ex9DBDj4XdoN/YfjERLUO7ATlLSJmn2dDDIFR8YgwEKE
i4EPmrpsy7BvJDTW5VXvB+Pv8fRBOgX455sladHQe0qclWk9ns+XYthtJ4ChZ9xziyYQuMHwVWds
THJhs7TwnLJz6ZXHLBIZUBZlaMxGDnai4MejESqzQWyfJQ/Vssq7GzQe/NJbPyoJmffiUG2QYTA9
Wg2/Rfa2ZyWW4TnWeC0X326ri0KqcagcrI7fyv8OkJU1o4X/pRggZd1Cmr55A0WnLCRuMr5EXzx9
uVWXLm/DW4hp7JapDqxDf0U04Kt2U3iLlQjTtBH+JVqORuY4OeOohn5Kp69fomLMCMFXP4jToGb/
YjIC9PwoRxCjTkQW/fD2hVbvgtyoOad+apth+MdYVUN8LVmvaI6rVLqpyGvsK3h7nc/RXoEWVPH5
sLYXGQ7ghkul34cLlOjSRPYHg0SV5dX1xKypUj+OqaBjeyCKHqhRjaWv8+XtVJKks3XQTVqqnqaM
iHou8vlrDjRUV+/s9zjIa4p1gbh/BrKlCFx6+ZdPBfRVJiHi4q2dM4He2c7K2ta6I/SjnJuSvi9M
FUAvBLoCSMo4cCumlgGcXHs/0gdy3tSbxw78j22t0pHIGNlMMWbL0qHS4zhx5WcNI+pr10mfqT2e
/gp35/BLae8ZJU04zQQn/ZAFfql32dGEkQV6/0fq8mh1dBHXhVaIlXh0l2eGkZCVgetcgOtjC+hO
0cVTlQ0lmMz7V6snUuFJIivSU9NmOWCJ1zBEOkfM5UOldDFaLsQ2v5Pt4bp9TEr2Q0cm96NitnPQ
RhUDCs4X+NrsRNZ4F06RHZpjQrNmjxiKcIu891SKuAZLrNIuG31CHcSMl4w/u7ZQ8vxLSHcY8d71
GogKwkAZ0mevE6d646YdxxJG4DbY6Iql8TSWk3aGbxqjSYRv6ScFbHxiis78eDmEsLHMPtIA4YQB
D7psoFMn3FAMkD6WlI7oUtGdlhA5QetXYjoAz080YsDC1YGkObl3BmBpgNwuyEMb5OrCKxMo8luF
3cD5Z5tnZkGoANnMoF2hTpJG5KMoG3L3OSNqsfIKXHH5jdRebLhdyJilh6ptMlTX5gdiDRqMY0U1
YomEsimb//rYHOX8o0Diyteuve1QVnj5dXES8ovmRKSOwXRLoWizDbs5kzyorZdPA7euPCa//Dwk
LCiIEnb8t9zPwnbsgY9ccSmzTx/X1Ko3eZYTSKZFLS8cj+MW/ZKacOL/eA8E4UKtCB97GILsC4b+
9WjN9OVzbiVmk6RejGAchCJAyDxjvJTTq0uARl1gQPpGfbv32tJjyRV0CsOm9rKUIczuM5+fc+Pg
JhjzDncJbCmpXB05Fy4jcG2wyTOU+5TqzfOJZb8+vuX9ts/iX0jsYsz0HO//rkvPyEphHFHJ3nZS
V6z8EfRFwmAhZR9diCD9C2fXlvAAoX49mGE7iQ4DJNVx6FsdMZcL/koBxK9GlPgcStbtJZh388kd
8sMYgUjSrKunI+xb3E3Ilh1BA5EQweZUuM297pdwmXRNcaLvwfH7FNImHDAmPTVQ5qKsWL/WfSWO
na+kxTiYZo1sAv76Hei0tZb0g+eKBlw7H8YowUspO3DWnZfrm8A0jZk1dr6R329XLPpPWHnIDPCJ
Wg906GBSV4mQZ2VqLwsNaUYDkO7JJEpuhQNEa0UhG/1jdvUupJRMUSxnLdz3EkzH4UUdauVQT7YU
RSbaFp7fac315JiBs2EQXazRfmIBmcAkB6OSNp0CyZfDhrbEfI7oVpL1z00QNIV9ID9h1yuZFqDU
aqCrkqjmyE3213B5YCNRyMH7TH0OQEbq7diNFLJxixO8AAkmaFFxZSuFSxDd44avb+1PP1YRf1hW
gbcF9bM0jem4FVXRIjIpyr6jkgKIPPr3u349tTPf0AvRlk8FC7utFoxGNzfKmJZsZz2w8paa63zS
MAnjLQxBPQMBTNUboDxpeC8FdkWQnhIngBWkNtF1eheCBYViviqVZGtBcvRGwMsbHKbidrPPdpo1
bEEKnrS7k9tEMj4rHfGjZmJlFSQsgTNOAjqvywdyKPo+7HY6OuLzG/lFfWmdis6IHqba91AZGMEq
02wldQi67shLeZK9a1Dxll1+o0eecgJVb+og4xF/3u+JKfzeyhfXzsXA7jfMgtSxpiBBiaEpuxHk
p+jiZcrlrdSNA5iqPSCoqdRc5Rj9pWK6KRZLISVWqJL7pzcYxgyoqVyoFNycDHaKAv5VL0u5j4pa
vSkGk/2npZFwsmO3lFoKVQMGotavysU5Kiq7N1t5ol0AU/sVwUUhxPzfpX+UMKOtXPj+Rl7gh6ET
IIpMmL8fQ8bBhKGTD7tlmBoDm3KDWTq/iN7F5DHPUATPl6fdNBzilJun4kiajvV3UAXWzQ07oUfa
es8khdPaZtdSKgapxkvSWtUr0J+AM7GgzvsE73mMtT5AyVDppQNXtlwalpnOvv4T4jM1a0P2Fnqo
tBE3VR9os9RKheq0x+qLigwfiKhCsn0Q8BX7thdCUakykf2abHSE5niTm8AABPea/irdHCm68Ie4
U/L4ms+Zh22D1dxZLF3vD4E5i6+ePxJzaL+jvrJYdf4mkESVDDqQUjFGQWAH1lMdNdI0M0lW6akh
hKHtCvIDPSV7W9tjLHqkYLAhmWyjIjSIeDWm9mFVs+FYR0W6NJ5WeeSVOgwbtH5M25lqeDWI4vJA
0DEbn1J8jhnATCuPr1qmL7ojTvIJhfZ8+G4vjD01kmcQfoWROSEF7rARMlusqIH9QLKoUuquhD1a
SlXFq0cDw0VsOTeh2i1c13mOrPdI+pxxIkK3S3eRBKGaTYa2t2bXBt4ad7K0NfvDLpohJPCMRgay
aJqbGRwsG0jJI69hKA/Fje1Mp6l/x1Rxky11+5jG3T2CcsIiY18SRIKUc1e4S66fZsxDUIc0lFZc
Knq49F4zsNoyMj5u6OcKeo9UNozfSrTuXzJL4ufT3IqtUgJin7dlXaJEMwyOr5jgzf7l/xIgNrZf
y2TdOtO3sNbQKBz5EOarbwOi2yh3We6DteFql6nACrn7xL+4QHbWUTB9IyfpHtGoaHHVmlS0Twnv
9YoTptLpOGUv/hCLhCiKPXLpc8m9tFXE9h+n0ohBcpmuwwuu5rJ/NFVMmMTTXNPPw0iR2M3c1TEh
j3uZ6S9XmTB6D1yUBw2vxLJ5L5fhVnp8GRtqfBWNNjiwm3WVQ5Bzy1hRxbwn0gXW9ophxCQ+cWM0
ir1NNM/nWLo+B9wvbWbh7nSAki3gTj9Nt5YCODN+W+5v/v/VQiNtG7DpM1qCw1qj3i+C7v8tSHj7
Ttm2NZqBcthnbP6YPd4d+6Q4wlw9qil6AjOXM9r3+6xBrx5OgcTI1uq8doCbQrGrZsCI5qBpbfVk
pVWZm9foNThpq87OxtsRGIUjBgwidmk+YlEEkgKba4pFaos0AWTvpyXcwukFPjFAa0k2GHrPBCSa
MK1NF7P9bDhSaAjMOsbFa/4trYlrwh0T+E024w5izx94qJVbfNYx2R1c54hvs19uGSIqsPKQtXbR
srm4vCkC6UbM6Do2pKX1wmV40vVhfmdweRVe3yivL1pVidZqPSZUY3xmyNhP/IZcOWkO+fk1ploX
uGxJdBQ0sH1p3z2goh7dAcu1Q3vbPL5tY19l0/DhC14gtGUYcWXyoE7mduJrrWAkzLZTKOXgPXKw
8GVFYXVG+nAaHW2whBT71FlBzJCp3jXu8AJgsHWBKo4EuzMHOJQZAZ0panFQJsenkJ0um7Y1FSQz
AKXADeOAxUgJd3F1lFYaDv++cF3V6wf3dsWZJeaNaCnGtasABByMHBmqZL97m+DdqwBfCUU5EcpE
BH3v4G9cB/0gOa6DUJJr8Bjh8IcfCaG9XM2Aw4k68azjAiszCVqQkT8eLBU9JkvsPfW3IBPeGUfO
0EJ7IbOCl4YNfP6t2ZbYL9L92nEkA5g3mX4zoB5vkrZUz4YL4gN1QCdL4joqnTrKSBKbbrv+v9KT
efmf1FAft0cRffDbmd21fh0ibRhI7NqNbZQz+imvnLpn4ftGLZSUtRGwQaHxTPEZhs4v8s2/9W3g
v97uri0KhsxSMd7DN8MCqHfTQmLpYBul6zSMmOkqP4O/WIr1HBD7HJb+OdpvtMJSlP1xMxDHETX9
rJH/8l09Po/TxzODBfa/mwtAMpWjYsrCqD3qGWWd7jkH5dekfoByr4711sNaL7DDHfpgv3wiUH4v
wUSZjNTFQ9CQ6uVN4HKOHWptAzM0SN5fAAPipJlGcloY/73vbE75fFVfy0FuFto9Xi2liEHe4VQY
NN+mFJCfU906Z9vQDsuvdYDTHsbLZDRP89Xt2bEmqpDu1hAt3+05IxiNbFSXnrCCRTCpMF2LwdcG
/rgx61HA3WSTJ6qTX6dRzi5FTy1VCOayx2o8uQi1JKYzTJn0DLDWsNW0IsORFpKIvU188pzhadkR
qx2NoVT6hvQGccfEZT2VbxfZLAzieBdcl8szgNtnV45aDtRWVF7Ckm/DHIYuYQvTWf7NlK2h9Uh7
dhMnuMpOYJnzucbiAN5F29ZEoWEmmpoc27E+yO20G513guECcsEj1/hmojzkMRbv3dePR532XQh/
qTnJKxU9/B7FUJrbYQFC4bJ3qDPWoVXPf8my4z1S1wNj3OjlZQC0hnp8FVrzqFAhPiCrRAK7p0c9
PSm/V0S64lWq2FkiRPvko67yLlq0osPReLXRsMO/ZE4g8pXFHIwtbdOMwgtgdhnHGspa5qqaZ2Mj
1SNsyFFvXQH5ST7qhdE6EKo8iuRxl5jkB93LFUieNjmJE4ReFip/R1naQIOweHdiCxoer0/Y5MOF
SrEjxvBE4KzKZk7P04erQjMvB84XizVUwMi87B5nN13U4pELoh7Mts7tmbD3ThA6di1lzeZvUJaN
soPzmVGwHGgML5Out7hXK6tAflg269C8q2CNIHwF6hwu5yqQBhFjncWBRZ29AlX4/yBEefifq/Tl
QQkuYLYVT7ByEVg7lXeEVUJpsgVbJaQ90UfE8ggPtzUA9Badq+O0CQXkDMmy9YtCxZXBXqXtvidn
0sG/fJV+jdRum/fuWo1h/0P7B/p7XWJymspIWq1/BaYvhWv1TK3j1NtXg8KZ+vg89ILVQhLmlFD6
xl3rn0O8ExNuqOenUfKgM313AraVV1pYQn6BJAxEvV9syxcOvajZbBQVjRm4yhmlnoqQX+3iVOgA
RuXaPKjinUvdYZad/UjTpqMxGeOL7ZgsZC11wweLAdY7RMI/jPxUnIvr7F4H3XJSaS1tJwnNozS8
dsfbT18IhWqFIaZdORUGw5pSRtbE01dJ0chcVhve4x+in5IuBml1V/pZC3X+rKc2PfPCZRiaPFuP
ckJgCue32UyHf3YciCm4I8X5GoI47XtegYlFd8eshdZCq2KQESYFB016t1XxmdxEwqtgE1HLzdGy
zaVf2jzzWa7eZv7+a8NJaiMw1ZxVZ+AR+0hjhxSxvuAU0DejBZXPkO69aJuzTbK+ZpwXf9kFieqS
WfUU4o4VpC9jtO7tqBT6Sw7Ru+bZRsqzkq5RoM2ODKgRuz+ZOOqXGyKGHJrUEfX3lVILLDQ8veAv
V/zWOkLCwNCtb1VI6/D2KS2JhTaS9uI91fCY0Q+hiAOUFUzNLh5on6cOTrNzNXd3JZ33nIN7Bcup
rH05er+azryTWI2CdQP6sHpvgGnV1ik0PYEY+cYBE7iE4YQaVIem0YJM5Cx9CzKCMYhSEMuQ3BWY
hAXC5MkNHYGu9VBQwxsGeyvQTs1qv8NSheax1HX7RZLqEedfXKT3MKW2iAjyg12bLFkwWfRYVvIf
7DNOsQQAYNQknoKUBwyiV8xVZC3ilzJIvknKtAubT7BvP1457ypXZLtqO0hURyMzeBlQ4+3UCzNg
78yOejQ70GMtk5jHianWLk7G/VIbZOCL3HWxIyYYJi8w4Vg0xjGPeViSRiAK/I5ZRGPRIldqMGG2
QXPF3aTxyk2+4b/4GVs7wjvjz9+Ey1dWTL3k1F7hWYoRVqzQ0ou8+VEdsnZMU9micG9SXYMPdr8G
/RY6Or+/tat1fCZ7Ptsuhrio/10rbburYJyOQr3WRn/yHUng6KFO0lo0GQyUsZe3+mHjw1sDgT+C
4O7bkgX/8o3KP5EVhPvN411KI/37DTLTbe4Mw/iGtwZ6wd4QUul9UY6RaNw0jVdJ1j2vf1bs+t8Y
AvsrZipwvfehDv2M0Uv/d0FvmFFaZZV80J4VTAjmKaUrfeJrJvvf4+KyU1BlZJ2DGLUajMh/sZhn
JdgdX9z+cxKRU1mCvmFEvrp9RebHvNQr+A+ZryvwiIH3tpIGhqwAHim8EDmSk9MGzn7Gnue16mbE
wwM2W8WlFKJE32z+qQO10wmio+9jqF0ZL26h/dhRFKsJ6nLCJ7ZMHB6KAl+Pm0gS5xTXzogUYUw1
HhMNZXppUnbAvn1A0DjiUnLmDpQdw0JoDxmRMP1mU39mvSWQYBW7z53OjCmYrADxk7MgMI81PgyB
s/UrFfFKgszJd3g+4Fv29fstMqm1xEc7Rm3qJk9F76nq9F11vFGh1BShhG9qdiO4+eQNYppxmmmc
F8x/fdUUrI9r34OIDRz4uX/LtY9S2lWEcTIlYpsjhDNUPKt/xhURUKRlS4/uenMJHy/efFis4Gbu
vf2ozU+wUqiaM3mKcIeARM8ndplbvc59fP8UYAHyFuzRWMbhiN3j65Q8Z47h9Rb0A3z2cEH1Smbz
8Mt6+vn7XG8qAaug4DaS63VwwjLkKNzt9dLRnJiBy71phOI/JIU/kbSZNFj6y0Sd4eFjBMn365vl
MVKtSzpm+kUe63cLhLyA8Hh1SL+tIkGt1P0Qllm+Qe05vC0x/v7ojTQAjmGHQOt8M/of/7f9wiZw
ZM7c80YxPbRFz8v58fGhhlyg+uR7Bn4TrPY8dxrKDMk+tUk/RYdsAFiKHzqHpGUw35EHUxlLchrC
47XBw+ZNo0xDRsjfim9O1WApEchDGLp758HpMNfWuOfSQuFUZG4lrGEz0ww1AyOeRdFS5jM/4F4j
mhliQfiGWoihNk1Dwm6wJ7lT+CLFyYXgEVqUWwVL9F6xvmRG9Un91dLY6DqpCh2vQN3EOcZ8owUW
AD/WsFQb3vE7+rLzgEviiAqe7PeU7TWiTtXCWpHbjKf8a8fZO6J6OxQJDGkaOc2gRJAFaH1P+Wu+
U8zCu9ncRtFuwbKASqQiBly1sqT8he5RSFuESxVRgNLKh+1tnHf9nKSdpA8zVtcuvhsBzxTCzCxk
ShBtbbogq9cjsMOOxwqvhs+NCUanG9AAfUm6NazGCTLEsmeuOfwdD/dhnkjuPssXKx56b62vNrFt
3c2vwb41rYhg9fHWd1iiuYffXnNmroG1yAUDMVbkk7w/MW7WXT+K+ZE2xh8S/fTC2OdUVeHUbkna
4pIvjfQp1OV9RMUTWvltcMbAgC3uZhLXO2Gym7/WE2SXJKJxtdSMPYvTHy1QuOQch76Yj8ivIxxm
fXdVG5YsErUoHqzpz+zLTfE1ZqQm4d0J4q4C7itCANwh7nsPo2xhq13TAiSNKnIAqJ3GUvgUN2Ne
o6Hw7Coq+BEykNIPdFO6uEtkZXckpCA3/LcRq5tgevam4EdYX5ay5EKiCR63l8XPNnF9N3lmI3lv
1gBsTQ3z2eQZ9sCdU95ErMigobp3NFn5RiZnrtBkO8orI+jJHSd3V2FaJXchMngagjWlBK0Vx7Jf
DSEvLNe6+H8pfuHPhRBkyqq1hu1bpLC6MBUwFc5N09lZFxyOGhOi+fWUQ2te/3gfiYv4AMUtxNLm
iRStwbW4eW0S9FX6vglpnmN1PP3kCukCLwmUetl1GjNcqdvswUF/YSdVjwQExkdyN0X6HQOXtOhX
JyIrB4QVMK21ynMEcDIn2Bi+MkoZII63wHE748d1ois8Ue8ErpMrqYPhD0cETq9uoylzNuNTcWjM
EsZ1Zll9PaWWeHhFgbr/hILTTg16QLJzopmE/YdRZ1/O04IvZdDDtN9qfYFiZ3jQwMbc6JGZHQVu
KbaWJf2sJ5AsgxwKNCxs48BBdP1Qmjls+I006GhPhTQFIIvW7MQ7g9jrPSPhIQHuW1MGTvQlZFsF
NUKlYIGxW4xFhUkOjoPXl0bJ5dNPk2aOnj1KyI797mPt6Pgzba7REiXdtFm/u23jf3BVRh1c5G3a
RICkxaB5Q6FBKaTAGhDFZ97XiNWilJIEu+iUXPP042KMHN0X8rdCHqZUHn4KcuvQhBBrO/nZGg+l
dDw+1P0dIgdBIvOo7x7SIcIDlRxakz+xzuD0d5BwHUqRhOkX57ZrIpcBhPhZNmGxjgLJkQidrQCN
aBVXFEDM9Py0BSUzLU+mCecWb/VPN7PyuuK4Ia9kxYtUw3fycZH9Ql1vCXFEePQqzQH+c4BU3IFg
SKoQK2N0Lo09BwLh79Pu3G7QxfuWVZzgjqsF8s7T8VjXf/SuwPjEOBwk8WfcYtFzhfe6ZkoeVLxc
OsjhoIwKUsrv1bj+yXS+tQoBvhCWEBDIy3LosDkmdX1GJKkmJgRkLEzk+t1mVX2IP0FHoWfb+M4f
iDspprXg+rgp/ILE+YMzHN08TlvgY53MYqTIdV+Xrypgkb160B2dBRndVG+2pC5mHqnziYJiXlOU
f/ZFJ3/CT3MmMhbyK1dI0n/rPQZqNkup/DId2ojEIlOYWjVNy1+LMtiHO0CmmjIy3Um8p1QeoJ7d
lC2f009SlywcMkkqhehUKEaWBLSWoPqePz7fT25e1KAaodk6lVVFfANVehBsQGT8SYiOkENzFuVX
8Tw9B0JrkDhMdK7TNvg6kGgd7iMuWCJqKYjkrvxrvD1gocm+lU/E4KbmSOWpeeTA0azvR+gIhyFj
1pSo3kA9kzT9Ulh9UCMlWTJbMC90IB3ttDeN+Md32V3WcyWLq0CqNouLAlPlYK0c2FJpexY/RYvM
p5G5FtyRo6mLMoni0VvpzFn+l8f1ytakRIp9AZEBVI2DOoJ6rjDUnYvy05e+kQr/Mb4lj1bZioLC
KlnHeA8QZFmnGFBkp+ezWvdmz6e1nRJ/uZGCJPHRCfK6P1IkSikAuniQsGWfxtBZNQe6PZDV+KZA
hOj/1AG//Z3n2c3fAsUt6gLkwUeffGcJilG2Fk2mdy1kSo2SpikT10fbnUf5+GRo1VSiYYSS1Zt9
xnBgdUFrLq9cc/M9F/1JPOzc0AbIc4wVq0L5lnhh7toiwK0hKIREZ8ysNpTF5zg1/vCg9wNtQr69
6vuqYLYkYGMO+A+ECxXnng4L3CQ1DXKShnlfeTv+jXRLmaHWjPJP/K+nhGA5Xdbaj7JVyh9Pjg9p
1HppYcNx4dZdtFMThMdTblZBRSRXaURhcqZsJ3crMhRjzJQWnt1qQXwOwEx7DK60cXvgg2XtCeBt
EfhsQ421kKpsfynYtq5jRbCRenf7KpmAFQa8DhFVmrjb5IAmbZCjAqv48eFI/H1Pg8UYuX6nN50K
cs4c8gcsPH5J5io/8HG63GfXLpVh4ssHBN0hxZyKY+4zzwZnYIrG33kCxJNrDu/JmirTorMqHjn8
f7jXJzSiDrXmVB6Y7zD8TNHlWhpqgD4513iZ1OsNxU6+bJXHTjh2SlSNVb2p2Q/Voo4r7luKBqMG
cAaaO3Zl8UORVY/Y1AqP39RrF8wCkjCF8j+mdNW+D0kv3KgYBiWYOpbS0zBzxiRzz1JO/rPa8py7
kL9IGCChHx7QuQlcFHuPNIJZTkMaLKRmzVKLPvGqIeTp7MLCDKDojOlysblTnOT82FVAyQkzXvBC
DwpBs4sGySpdIoFmE0zpoCqA1eGbeSbXw6QqQh3IYVh0FwwGfrw9W2cNaGJxwzWsFIzQGPug5+7H
JglSOrMhL2MSF3p94mvZLuaTLPgPwmmHRUppEroVbIL8RYj58bxoNYD/yvnl2gLNUQWDE4tcc1+4
xYW4nFPGlTiiXsgXmSV17ekGHyZoNke2qGaaBSTvXfJD4Kd49APkHM1h6u/1w5hJWrnAEU9lPE34
yd3hrjhVe6tjMpo+bKZXVr4+vrZYR05iwd1DzqLb1FKb1i4kySB2I+EVF8R2x1VfZABTGvwTK7Ve
LXEbdHuAjNKlxeJL8zihO6trCPONXWdHGrZhxkzElEoHSKlaMs1JAlWIFNCVZBXbuoQg3wTcCwNz
zqbAL8qIAaW86elj63YBtmQm5wvXlnFQbY1XswOPXt9PegNSIPA4c4/JifJXJljI3QxmieJ9/Mm9
swX2LkyMqRl7CznCidgdvmZGU/0nSEz6Owsfp9rdS+yZbLg93qmxMZZlabWCTzuNQOClXO1HqiGW
IwjfxSl2dpg9e1zmTj2WWP91kWjNpygclXtyn7cBxl6/mDEw6qcqsnd7Or9+ngQk/VPh1My0yCZl
zSQhrKqYEJJE5iHdSjtE4Ty+OuDI+MLeaHO6qH0MDaTz6xsKiJ9mX+8JT7nyHvd6LT747l78oWpS
nw5fz5nmw9dH9bHTC4O36CcAKW6/O+sgJomLiSG6LasRmtn4twqhqu0tgAy436obswJ5xqyMPX8I
Ck8QKdFaA7Z56SIlGFX9GR771s9v3SqW6byO+l3vTfX8y3KwwXne6Y2NqI+ZZAhf5Zap5kVnebXp
JQts+jOHza7kQ3GQe3STRl/ygOBdBLeAmdv7+4vTsbRbeopUBjGAn89GPd5+Yj+G8mK7SwnJ628E
MOaXL8oBKnEI1mlmPEqK3hIQZDk3qU+6GMp9kK2xt8tPslogABNa35cqIK3LvlpTF70RCv0XFC4y
dGSYmCERDTGF20CJeh6WCm2YC5sVQID4l7GvF3N7TfWZNAk2ArbIlMs3/GsfxK1f1Oe3Lr+TZ6wq
1Cc3PUG46CWllL45ZX4o7Nvcm2hIt2f2eOjJyh+G/9oq6IuwhdP9TDNF8Qu3klI3Fm9Dikh1Z07A
CKuIdckCqKUhQUjYy7dEmR2iv58Uezc9MLw0lK6uJ/BM9extNSjKg7pc2jxjur8j+PcAivqAs4Cn
oXxakLhsqau3FLCd5NpYJILxIwc5Pb4fM4IN79x+RmpIzPvyXC/1/Uz63ZG29ERAe5Q9bGCIDvhf
UOLlZ64Dsk1/ameZrZg0eqGVb0kwYqJ24svPFOzaa1Oz/nzAASGYk7B7NwwaGEHTkjn/FwX757XV
VZkFyb5GlKYzJ58+fA8tiRocIH4NSGD1Gvz0/c+bqkQfRzicu1KMsihU9/Tx/viuTFZV6KvJVNf5
aZsTmQDRegYhJ6ogq01wxr3m2TOH6R5QjqPl6WIlvOsbbuJChatqfr8Ynfhckg5v75w618kGzTx6
djdHPTue3ik/F/5pPXJF0tGyO1FgjODG/Z51AuFcLSBV0dMsv8aQ4f902GRKyE4Uu2vXCUPOhWha
n0v+fOcOml39bhbnw25ATE7Erhk8fathvw2mdq26ys2VgjzQEB2DM5lNeWvx5oc+cFf/dQ1xgiF5
+O6XHqr3nCuLvxIY9ntsY/muaGfRSzIV0YX28Ihzv4BJQT7g7yufbdH6p8izM3yAMp8O+HzND9+3
60Ts/qUR4jpEW2Cg9BFAnSv4fCn++AekNtm33kP1OFehK95BrLQInG2XYL0FExrtBTxi+1F4sG7P
X2IZAljiYEs7Pf7k3Hatamn5xChTjhdpFbXqWyVaE5Pg6P7wdXQ3ahqA4wxXPn1qtQx74cQGDsLf
U6SwqSffI8IHLm0qHQ0OSuMR5RcSX9t2GvV1W2700jrFaw86DPlx+kattrVxEMG5fA6Utq3DS754
z3nZ/+Piq0pEXe+OJBaQTWrxE0/J3E2lyen/CDIk28RlGTL1mucQHOkOKM9yXWfHDDrghJ1radEO
R+y+lPkOhWIQAUnNGGZSdEdHg7W4/CsX27MSnhDAWMiNH9kcXUNg31nxLYI9wnWc9TJAF8FTxZQ3
HZJ1HbVtVqwZHBQgR4lwuEdWwq/CJOQ9s+S5hFxQsct8EJGJPWr4KnFysPaVoeqBiL1IDxNAKweb
KSvtcT8yClUh4YRPc6euQiHdBhrKN2tOmJvRzqwCgNmULX7Vx0LRnXgDxTl6MTTeB83qgZXJaiy5
RzkKNlpoaJuS62DTl17jh8Y8Es+otvQVtJQKSRofmGfhf+BtywjDfanCVzenoazljTmFUD2hFMc1
U4uny+Q1Oc+TlX5Pr08PjxGVPl+9rKQJG3Laz07pJJZCuziL+BWOOs6MOticUwfBvw0cnFeEyVVE
5C0yU9dB0NZcn/52OaBDPs3lSQHTEMslTaT18idQGxNtFbd3uFrkqVeHJbBuTWH7Tm83V6SAt3AB
LabUyEa7iXIq5xike910XKZ6tdaK0aGy1FedC3UiJZ+qN6em1T2/xrRbySmnMR5nVrx8nJ0i540W
hGDuptbHX8IvzpoOzPw8AcuTGWDmug5UXq3WYlTfvwfrRP8hd0BIEiNoYtU1ghYa+yUsxzFnofV7
S/CYka7Me050Vlpp4T70As2K03aczKc66jiWkBe18eDYCyph7yGqFfP44qqxbRE38aC7sqs/uA2H
myyIbCvVgmHtXzyEZWCbnBBmo/NCdGOT55ooL84V1k1ApPxaxo5l7BvSfllL36W46e3HyPb23yOO
wf6+w9Qdq6bjFXNZ/QQnT+APrXZfhB6kVt0gxusf4oyD3Mt1LDuSicwfTKWYNM6CUNZ2Ok+zr8DJ
pgSAgEsp3icQwVQ6/rmOFMwVvIXEEQfmB3tX7C+prDU6z11aeXdu6rePc3f5iwBlwt7YkBN/fqzR
7HBL6rvtHmCR8kQ9pStkLfk947obMr0uHEaYa34oXArO9K7zgxoE3IyE0XFJrmQoKsdSy5GxNyH3
+roGdWzmgU5Zyrr79QG29MEXEW7N0am+2Q2lBTaW2lF9cX7zeOPiVn6KojKqZfgPQ2HrOjt/GLlO
p05MW3WTYYQQ0lkQ3zL2Jm5+RGlqXrs/JU4HTI5cp+nMgQLt+4xeHVYG78Ff1KLzaRy5+txaVois
eGcpcUQt2Ci5qBMkbmmXKhVLzERngSx9fBdezE3A+ICl7/K9iWILdAPQKgIFx5Xtkrv42tufzJLt
J4ePMg7SptD6jy3LUGtjn9LZM6I88zGS9qZkQwJvAEqwbEKEVOQ5gi21xlmHPvVOTY6jveNL6t6x
gJuTFdlHis0NApdk2+uIO3XU9pY5sbYiZqWNbim2Oadr7fsxv+YwZsZ8MmZOl1RVFEeADrqBRi4F
Dm3xdBhKLrNd4zcu83Jk8mwoDGqC+iNxf2gTKflZSPLVb9vFR6btcBgEyD2GlQqrn3Oc8uzk4w92
72JMNpyCmWPyu4sP2UI2WuqgyjINpS8q/Ol/S17ZTI62lNbk1v8EFytAQecXL1EgipU4VkRvMiqn
kC8flIE5VlnhhEK8Y0h/UBfDNfUT5UInScH5bHDra9s7uW9pAAK6hU90Fr5ZBEPjwqv2u+UbUwwC
f5nqzB7eyA1j9YKVloIs5mPEh4nnTIcF/MGZ49s9p0XT5mEjOMMmGvMu7CZDnYtFu8/a+o3FPw3I
pkEKteEr7UD83/RrTI4UwKEu5H4d9f0adzhJLms8QrRBsVzyNG2dIKcTiHF12x/2joEUJAF2FZZA
7Coyi5QKLksWonvII0dVW6H2G1PF+fntwLZC6lZGy1aOqI2dV4eYHLSFdkJkekl+nCWURkLyMUoX
P2G9+dSYhuRBHAN4tffBx0lp7m428yC0KN4NsXoKAsapwbnymLHY0fX89PuTJRKo6sHserqJHA+V
KPK5T8bcMa4aSCPc4cCQGDDp22e0uhyfv7bA7E0OuYeWFVu7xomja/2kZkY4ua02QEI3WHs/02AS
/itVSXRmCG3fk67vclEjuhBiaHkBkbER3bwNaRhjyvzlrsqT1sw1pGnJIWe86MGHlVmcVuNYKLbF
tn7T/JWpTldXeRQuotPaB1DsmL7B73Lo5MhCtO+rhUElrxkIvg/a7/Bxrch3bLVUO00KWvaFmc7w
0J9glB4tyF6rpE/trngS802HWBAHMVF0hv9hso+S/vjB43mbNRaCBdBsDn5x7rXiH+Ts4un8LnNS
UhiDUYoUTk1FXTC97MELwA6L3XaeNkAVtf0mzjlxTQrHIPq12055SEFK+dl2vgsUyyYFMsm4RO8F
ZUOlL1G3s0L7whHfEwnKCRpBONXmOEuTi7EaUqeZWIJPHR2ajVJPouKp/2aY7U8o3tcexmkCBQQB
hou6h4NBXSEc4SK7J/nBa+Ccf9f0oTiuWHxx11CR2fgDQcwl/mDRTlaX5S1Lis/nG57qwF8dI+hx
6Kvz3Z5K1qx44eCqJxuFW5cq9/yzHUWKbLAFf09mNXY2+GOe/QHjlDdbQdE1/uGsphqulpkRlvyx
vxYqqtJa3cPu5VhFzrQ1DAQYz5kqp2nVcDPN9TWFZ3sYTlXKvgSwOKPljrQ4228XmNknrV8JI/Fz
Tde8a+Ee8vtZKqNrOIs5hvqZLijNVHDy44NVWkknbYP2YGscfNqkmELD6pFlvWocYUsYWW6CRIGY
IUE8UeQG18q+IDX0E+492gY8r8i6iijIQ1JIBMcNQCK+kK4yvbezU9hpJps7E3zKcvwgB3wU62m0
KCQE8oIVHHMWHbeA2jck3jWUJamMDSM3f46Hy8QwwZACMvOrHKwZDYFjRri2xUFslMEGS5XBZdIV
pRyIs4vn9iVF5vpb8Bf9BlQAsZoJ313Ctkrx8FLw5nWsjO2XllSRhu8bVlmqr8lQjHSqfpXl/Sa0
FhafayxnDlUbyFJWIuOH4/UD7R2X27BoJrvovwDDUAlCZFNghhIyg6TQE6Hp2pFLZsZgJDSJI0ir
PYNcyvI/AqvzrflqQKq1sOTPYd6Dxx90qcECdJ28csDvMLPxb7UwPlN3amYk+JfQ0bbWhn6cXw6L
pzKc5zku7e2ikDRfxcdBZMKb/kh7PZoWNSEW7RRkT90AD5c89lAlbh0MQtFzbsaMwqjgwh/vAw7q
n7soE1p4/nuc4T6D2wP4KQZBPZOCXLzygnP9qtHH3wZzBXhCglsTaSzLe9gzw/SuRDMiUG1FTcH2
dpr5T1A72aBZyRFmWaopAI1ZnSoRbLVLrWUv5OeABW0JgBZDa7jeuMojXn0/o0mTDaBVRZnZt6gy
5snu0lJSp+xz8413vm4LaFk2liwE8gezjTo9h1YSsq6+RtuY3/3dE5NFdieH6G9v09MlRbESIPUi
h8jc+ycMhHNjh43L+n/8wzg9V4llyTQiYZvj71+/INrH3+x4N/Mx0/o5ERd+6pFba/ZePiBGUbFd
61f9E8n0dwadZ6uvn8r3p/ayFk3SBvjN4KovMyote2IKvXjwgtzdsZ/tR8KkZzW1u/UD/12oxyB7
CRpCeVh+vMnk0HFuXR0OWbR8jhUlX+OkvGhp7Bj3QmC8Ua1m7EE2SIahttICWPpiTsX07Q87uJ7Q
bQ+u7nHSgWPXKusgWOqXOEkSi8pg0p0Ja6dpStCVvJbsRKL2y1KLdd4rbLxhSqL8Eh0HJbHEvjIt
AvO6qYSsTdNNMnyAtGQG7qpobaNfK653/1/EsADoX8CpGEDln5dhfMdsnwSooX+uZCjwCbFWQn+g
hetHlfCS8ACYr9iPEERWsZm/62mtzqwFt2HS2Tv1OLlR1mvDnuY3kHHwaam/R5E/w0XNfJNSmtWj
qi8sgTRbDNOr+PDZi57SQkRAnOFjsjR79PQjrwQZ/uZ5cywBBZjmFTb7ZRfpVrw0ecPvjuN/i4CA
z3+WGUVp0Sy81OSZ8hgNida6mDQ1xDPJFERTwQFMTr0icTPqnO4cfhHouDvc/Bf0cPFnD6ZfpT3w
mm0mDSzrchFCI+F9h4SiwvJ1Pk6/BL76+P+mPwj92uQHgCiHCzb+i0Ug7qYP1yFINAQEKHbFcjWA
WJMTssCI55oXOJjsZ6pNkTyUCSFa8zrCvT6pXZFK2z0Ule75yaFrLtsFcHx9Fp0ypqMAbW1AkyGw
LtCox9YS2hArirFsOjXcKyc5CllltzLJfQQPfSQkphprYDuOGD82qaE7/4x0jB3uBnWsvo8Yhy+1
0bCS+KajL5gVA1Wjbpor6vj++6g985tx4zBkmMxjY8t+TG832Q0kfLKFmIF9fxsRqKTlzQeWr6tJ
VMB3q4jY92Ry2VDwCXwnE22VfjtsR1Rakp8+Do2JKzhz8F5VC7Su6O5EJuKwQy34IWu9oWtrdGFD
FxlipQULiKXOOCeO2cee42a9eiKUNVvy0xDa583ePWHE7rKr3aRtEanoNmoskTuu5RAaVreys1kq
XEKlux3+Bqfczb0+CFBSnvO19NZ4laUnNwWtOyB0nQEjmt52IUUhnnUpAYiYdE47NpsrcnS8KZFR
t7nh9ftyc+QuoMq8CmiEGNjUomu4Et9XeKVjZVrn/qC5zxgiHa2TJhBwbo56AyxEiz6UQPs4ti01
296VJsA4R+DsrNZxMCb66fnvp27oNMx7p3jL46IsJutrMdLCtKuhcZ13uN8oh68EXVx0EkrEjh5x
UOElQbuTk9DlXbcXQEQop6kTA5aQ/M60ZVfZo1RxeMziFludi7RUKViVN2QuMAPdolR4U9j+U087
oiCIrwBxw+6oj3XsX9IGFJOw+LyyBa9lQJgicUtg4Ft10JPXYcJxiBv/e7hffsYucmDGNxCqDG8+
7e4jMg9IZHXRuGsHIjQ1ehe63DmFxu3F24Mzh4Wm3zx4Uh+Qh0OILOocnWhM4lDymWwBn2LKeaca
Yn1pNqijuYh2KPGh1N3wdesJ5l/fR7KvLBq3MtHhVlmgcpUozM5NhagitIciD4zWU5VuSrUrcvt+
97U+ajwfW822sySdZdSui6cjbf7ko/X4Xgl0YhE3+1clSL9KDUM941BlAnM7HSCYehkX7qk15DP+
DilomXQqCmDDQNSo20v2ZVIYFhrFTM5HatvgahaOTCvrTNS13q+lTkArqVi+dnmIe5AIfONtIHqN
Km5c9K24JviUPiJIsTypMGA8GZ01004cIRWbPTfIp7o01L3PjsUYPYg8A3oST3HLpQT/WNs/V7FR
Qu6q4ljeyKhQy2Dq3IFiKVG0RaprsppFeAcYERuPUPK90IXL1992qZpb1XFbfo501Dqi0xDNadRe
En/KSGIzAx/eMyXWNyxq4H+IiCmZSbkOcrDAdqYsXoFCHZIow3AqCkIM1Tpvcbt3m7jo+PehmS1z
Npa2OVJVx0phDiKN8NH4SKBf1x4QtTXamUILWXVXn74BMH86MqRKJRaHu4YCPfmQCPpkqaRVapBu
FwCpIViH45fik0iKLav/RrAelbE5dxcjaVABAyc1KdUarNxY0UfIIPHgrfzHVXvo/he2kXfj4QUl
1SNtcIzjkebIq67LiQQdFnDzdoiLjtVqqIkuwuzCJ8n2uWLoilg6Mq2DowRNQt4yvqbxKO9TleGk
4qPpHQf8rJhhJXCvPJ0Y4rNEkMSb5FvrJBdc2gB9QkbK0lYkBpuV0gZo0ju7hG3QwMaLIhV1CnKP
EY2dql9PmfELB0+JxlujL2vA8SDaegxeMedVTtq3ZbR9E77rT3xUC62hv1WhVF+vZnpEy2A06/gM
tXHgXzBSl37dbEAUK36T7o9sagUgixyZgqWTp1e+eN4/KjYwVpcM+A5bChhgcWhSieg4rHdksMZ1
wRrWP/bpX8L/91mjR1M2JcNbHg8+iLoc0tq7Vni8v3blOufqZrwvXyZt2b7WVd33FUfAp6ea7mU8
9HnzVgpIoGMLtU/oT/DNpyIObRo9r+wJO7uTxF0sFwvLTQAv5S3UzmsBE55ZC+zFthll84iFh8pz
Qr0ZF1nrxqN8LxDuLJ9vsFMf9vxAWFFLPDcLNyMha7FWcMNC9TEl+2aMlMa7JxwnxrWUGnRmoAHB
pJpQKEJDzVIKyDMfYzU4DPu18OWdMK+6sB1LhVBEG0YTcANhTq11LnCl/tp+f7pxOTi8wNvA+dba
p8+TcrA3a9LHT+y2D6fJ8j7Kt141K/zj9t9ec9T9E8WcOS/kGw38XRbi8XkDooMOzQ5L+VR8g+/v
u/iZnCtXZahCo6hLB1agoHmYhlPI1ZYW5I4F3UcYHNtodFa1fYvk7+TIfZDKjUA/dWw4f/j5Ukw9
8g6dkdTWNbdnboTTt2NIoPUm1oVue5qPPJbQAKOpm7twLLzzIFfZdvwy551biSpjoBFU6O3Bn5Lu
jXBVl/1etR7fZeU7RFhYs5eEsKo949ZlvwRJ8Qde8MUeUEhZLdkleiqFqehL2SP2/qxBMa77TJM5
BJ9ROuogUBq5p5cOWTl/Tah+W8+YVupaSMsTFI3DONIkjUzuBnd12sqEAJCl0GYqtLuT+irRV7GG
A2pjYfTvBtGSS7QkfQ/yUeo4iIL0owLTrsxaK3gNC5LSAbHBkR24GG25Nut6wTwofXMG/fflXTwr
3h/zyb5GK9JhycnZ7TdlsAMWKwDcQyVEW9pzl/Q6DmhaGDp5sLbu/JeQ3rZmly4qJ8vaZ/AtGTKE
Nrt1KzzCJuHsDBlInWsgpa6KjJ2Z6MQ7Ax9akY51KuDEJgkXfjJRYlbjX31MwnHJ7tUUtOinRDdk
CeZ2MFXUNdBVdAftTGsxn0yeiJ5ADIM8xend+SVML5xPyOM/5KWZqQQICGWSlGkuaPrwVa/W/zGk
q+fEUg66c8MIWVDTTBlrFdKjhk87NjXHsVVnr0mJE58NkfybXCekgq/pO0Wfn6sRi0QqJWyyuhWl
j8P02kJ/YWtTHia6PF6Q/U74XG4vjR9o7vvpyA5QOboxEMEl+ITxnzWR8Zmm9ZzkuGA08p9V8CxK
Z41bcqDIv7YUyvLd2wd9og4OyfdCdbynRTkCLvH1Tdoyp1OTYtELhHNYVY7zmKa/cjef5+LmK10w
CUbjaeQT8P8Vzp77xrNVHz/PifmbDbo0BgnQzC1vepwsktlmK8ghs535v0EPaVBUmB8mRjdyXs5G
aCFatJpJpreMsL4AoKpLMLOL8xZIbhQP5EcS0JT3nD48JzJ5oPTE8PMJ1U584JojVp4A/dXdrCcB
EWvYmDANsHQI68zjaHjfeJktWpl/RgQggRz15UR6+M1ECOP+/o4Ag9YyMts/Ctj2i9/a28Vf+EtC
9GqT0TSyWODkyhtBHZIQ63tlbznxTjSPCoNGnRTM0KnxDDbLZu2v3p5zoMQDZHNOc43Mi0vDXXV/
f+vDbaPa05qiuoQnr4GfwuR5Wr6IKbEj+fs8hwO7R2Okid7c3bNHR4mji3PoGHyL1S15qbmBvEKF
KAQA9BOdYGnqqHLLIhAaFjoFuOga8n40Yq+067MdWrDT+pYAnYEzriUBmAgZNgNTD78tzYw5pbQu
mMXLNhTIOiQYXTojyOEEZAJ1kvM2jTCXMS10J64FAslBPALrjSuQZ6axeaBORRjTMqob6HYqqpyD
WbokcOlgFluYnGOoGribwWwGQTmTVM2oB0kpX36lguOArE02wk+bQcXUb2Dq46rkufh89v2JReZ8
HRhRxtg3EpItGE4FvUQ+fXgxMDMVU+jMfnUzlUoJ1qqcHWusS3WmZG3xjiDqg5Dp/x9pDAyx8oil
PlIjv+/QQQl4bLBmfBt+QBfpNj9c+yw5pU4AOxLYR+yYv8eCL/O+LOicJGIP/tRLR6QDmYSNF8iv
4O0ZBHKmo8EUfvrcD2Ej8B3wj3bnu44sBCot1whSlLa0/WRO/SPIFrOhXiaLGGXfnO4zHLR6zgxM
fysHYbmqI0pQGrMMpw+zO9We87uVFt/bIq3s/DYixbCoiOHLncYNngLQYtmaHp2sIqNj9dtrJS5S
yCV/5FhQEm6xeEOY5+lYDNeV/V6PZH22TFmgyVqOs70uRiyNvPOEbi5WuHAkyqfK9VgkXKRUKNfw
rtESX0D/KlvRU6SCwjsij6K0+OdzKVmrGyrhnVi9eMzj2ubkfFD0g18Dj4FF4d7oW82WwhWHnZTf
gPwUGIbWTnA8e2BSxnoeTaBaL1lHrBEKAWjpkOF7lfh0OIgVXqRHopFrwao4/Dmh5cMOV/4oHXzA
p+VFrMdQK5bZEEIag8IIRqjGXaioBw5i3doJygVseZZFJ+RyGv5V9jdduSEUEVXAE/xJx+Du/mIZ
pTzv54TD4O8ORf6lD5Puuaks8AffOCzhDSjnTmIwuY89pXUvonm9UvEqC+GZyKQV86L9oItyA58Q
ONvGa/3EvlFBUiNdYb22u9Zc0l561AJq3wxyxtlhtrh7v1Qn04OdJ8OtJeupdsma80hCvKrj5OWR
mdwA9O7ddbfNpVgN+3Xdv8hGp0nhoPAxvpMKFGOzSsFhHJipcR/0Ey4sQxXdi8xzgUYYicqchESw
KivTDRsAq5Yeo6pGIrFvmTtwu+GdjMchyqQ8swL8/NplFmJVFVmR0TN8GGLzB0hKhmnPeM4jKalz
kfPQwZN3mv6Fk1qdvxGn5ZHAzil8vCL+pQqjcFw+Nl3/WbcQ/L5RsyZAERmGBZsoRzX1U8Ycvy6H
1ZYbPlO+9ygeVJ0YCOJyIl14X/KuMCtjQ/2UiOtrp3YJGRlNsmUyGabmWqko7PWq/wHHC8BMD5vR
0XunbO8kBw9Wg45/5+hv/DVbBKlZTzgxYeyHzVpiv+ZOZF3//ZP99ddtG42wOCR71qY8nqdKcGwB
Scg3ivhrlhSfoKvN8K2YxrdYuShZYvAjRp+WDD+wkuPvxNs4peNsj27YFx0jeQw2PdZHDyC9r7i5
ddLQMWK4JR3FAvAsQ35MAbQEjaeIiRygq3sbmCBCGdWfAtS09pwJWAiCLe6lTWvzHNPPylWFDsQF
bXveXlV5Xw7/1jeBSLt1bNaJ3M3/BGn6Y1uZsOb+CNm40wOXJ6Jqhv6wHVuMySrnj9dfzKuSkGhY
GHbZFwQPTjODBtRD/DnLLsH4zaxOuJe7tgS81WzldHLX6fVfmB1DSOurlLsGYRbi6cbja2oTMDT9
2WIjmYjdarV5ObyNNTPfSqk1FmeiUpKDxcIqZo1O1Za8HdtQXaj/0uvuhEfpl7Jpw5WvV86tVihI
m9ZsAlxzo8sIK+wM8lp5a4lV7ECUxdukpG3jIhalMBEGiKGyxkp7wfwvZUPyKlAuMyYOTcD2NCVa
8KzZcrOk/0xN5+4T8zmWFTATb49aDbewIN3JEqNZ6s6XPEqQBY/ElkOv4FF2z3L3F46RcWQ9uH1Z
r0RIwZ0GIpfS405GwEdySPGyaDh7LUZSFKffCRkg9VaURne+UL5nCKtGnEz7/lCf5r/iVVxceFin
2RXs96i26mFV673zM8ZWyiPd1m+A9CQrRxvSKlZoiQdnS491H/6RiiyBzYNN+La39PIcsuCYJFr5
AW/Sz2YvCwZGf64B6Ym2gOfgELNo0MTmUUYs5L7fqcWyOA8c/n9jYBmEXC/Tk3ZWXwVdr2yN/GBg
L5pdtwSMn8PUdEPaBrUBK3s6DUvfPetYlKL6CnUSmwJLDLQTaz5m7IA4KLXp4fW+Cp+53jsTUI20
Ga+2b/ruvtQTRSKRIUQZB29Ksz8r2ljzCKBz3kPws80Ij55MW0/l2zDMs0IBsVt4kO7rGOyPM0b5
j7tKOekE9GpNjcc10Gwo9ith+xSrAGtgoUIO8eTKBbWorEzeRPPcB/wLqPjPXt2cS11GWksZlZT6
vNd5x//1Pmo4oUVal+4AElp+zOPWAaVLUvr4nrnD8ZSIsbvOuhZkTylAdCgImmf0u4FlK32aGB5a
zK3kXU8ge/DrKXXZJrNWcCqW6J67lEHr6A81MpJAArLngCfs2B60yLjPbOdVQOMv7vcMa30pHGs1
ux2v3iYvtfLi98QMKtWMbyO6dcr82dIFvDSaJ/Hm8VnY9Y/sk6X+55CZjQS19RnPo5hOBb73mr9Q
G4RNNBj8lT/WYuEe+6JIfwPbP/vMTqXg1zc68Yw9vVz7tSwH24BuuKvR/RqRgd0p3uHhzcZ5y7Bu
rFE0c0Zitv1DG/SAGFdNeLqbok2w49nfXxAdKaP4LjJchD0qTgrK+GHc8w+dEezH4QLRuvPIZQ3v
bbOYqFMwh1iuchuUNXwy3mlY3rFkH1d5c8b4+c/MHTnXDqmn/tR88N0rGEC5b8qsSdkJD9rnyyII
eM0qJJR1k8/liOzh7Xm+W/TjP3HnHiERfbTgxVpsBHTKxLKFSYKzNtyWvcHDgBfVcaUMM3nFRrT7
V2IKufcIbgTV1uz7FqfyrCuzJEcIjTqvNXAFw0etTbK+8KQ5ac9dih9v4c9wtOcz7o+XthWPgTdf
54sGH3D8ZugHkXRQ4crLR2loFauMW6Jm8DR20AAFDuTQHRJsi/fAHVS16QK1OK7yEuUfbQKQxfch
7KC8LkRiN5koEw1xBMoBC5GYl460BuGSY3wdf6lBaSp0AluqrlQN5LmkFwyx87ur+V+X6c0+bA1V
X04Bq/ct7SZpbJ05C2ByrtqlptO0wCri97tmpBRoumig7Q63Imb/RiLloCdpuEacmj1zNAhIeZdx
gg3geGhJgXyVT7TaxAkHqxhoUMmLT/gdtQTNqPBaoPeABu7qN3fxXisjcPTHR1gUf+tcSchuqr/H
BQQI8uIw9H0GS4Nem/OWSxdTlMFx6+Nt9KO0DBf/7Xdc1UH7eC+S98QWFOIhZYHrffRR9h2zPo6g
JKznkL1ExjH4CQqO7I9dSnztRdN15xncMO35zK5Rynfjd5iNo8pAhcZpocL4OiuLgaBAg5iWmcQS
QtHzY5D9Pu1Te6/j+Rq8EkIJJjfcYES5C2cY/pl/dB0L0u18pIbU3Or5TBaOgomQ3jDc+FzWxoN7
vB0dsfK3BtRXibFAdUSNYZgjyANCB/Ahc9dUc30cJrgy0fLT30wmT8ez2AW/bdNg9yz0pVf0gYMz
7p8VHbj75hI48vGB3DaPVuJF4m2JHBiAGSvNebEcaosRwPZn6GbNfds1Bq+Wv8BW7DLd4rkoTeNr
7sSAWTqbklGApLS0wo698X/VZsVVJHDvObPb35qF8LmFQbo7X1pOyTHv36qyeaX2jgv/t0cJt+qw
9d9lo5VXdQprQjysDpw/9gD9zlTcm3Im5O9S7q9wAekV3o81lZbu06/LXX3NqA9L7V76GXGXNs5v
De3sidO4/UOONNRPcdja4QV1U/to9DbgjUe/B6TvZhdeOvEqHYTkA7VRtT8C395jyBZf5mMzX0Qr
7xFgep2OWF2BGcTq8+i7ugfH+wCDW6FRuT50NWWsD70L6Wt1wgZUyX6igSWIaA6tYZGZAsj+2U3m
kQEH8yaxlmZbhlomJhhMqN7q1K9mLO2zNWn2jyYNi74Hdg6vfF1fpGDEeED5NhHhqQ2LefpU0/LZ
gGVf3FnduDDUCrH6s2YplCJLPPVqmAGr+YqjUCFQk4NbMW5QzZg7jPOEg2DkboWvZTGYLZy7kIzY
842ETRbO7FXL8P3EeREuOYPbZBxriZEv1xFV2gX2k6Q+DW/GrwYYl42h1nf8OIyQPjmReOIisvou
eeauw6XFOIEKQ3/ttfNzBysiPXdCvFe+vZEfJpgrFGjcgngggLMolfsBvHeTvyu9U711TrXzuVq+
hy5ANuiv5SLaj+dKVL3ZhgfwjdUD7doFlweuAWtyLJsDRMZIdNnWSb2vAl6rjtouDFhVxP1uG9db
c8rn6oFjfb4MPQ+ntJRbPsfvQsO0qlGTQknyTXn10QKnhogE64cjLVmPNUYo/V4QqVZEZgCYgX3t
Pk5+tKcX8H3Xt4zA+SA8wKJ1RM1kD1X9uKAQaZDpuMEdCmy7laflUNbgh0HS9i3L7UhQDKN4KCKx
BR9yVhr9UepD2R10B2spVc1ct8gcwyU5ccokZWOQgAFBPgRe+Zo46rG3dksvPoazqn4W4vsUFqpV
m5Hv3/9oMB5zNryio4Gqrz1MIw0SkurMyZRmhEt+bEBGNmPTON/rWNFlV+zljQgB4XLj/6PriySM
jon0norKztZzWd85LRUjyALRbgOaaB74S5D+oivVm2L7XcB99KmDWEKFhacv8bLLThPginQM0GC9
JOSueKOPsHj/EEV3KMdUXwXvbDVslH5eDt7ObMEIXNKs1GMioFi52Qwb7emD3qo3ssP+lZSugFyQ
H1PwE8Kucy5CYFIC1WthZnJKFA1mT4UFtIdtLZ6R+7lgOvR/ygVzZG0f/1EkWyXz6gb+RXcGjVg6
sZONaMmjCCyVx1eSKO/q1dLu3E1oNM7p62tp67unWphg7q/qZn5CTCnRNZKK8LHtU8AG9d/aP8tS
KC2cRiotAH1YibtbfqgL+ag2twM1pMalzlsKzhnjCY2ynrk3wy8oR8E2SVf8TtRuAIEfZf5E3AHg
Zh5n8IkNDigEcTme7XjbVr5MVqDPKcHJloaR80Xw0cV84jkZEznpCEm9fEO443DkaP3+5KKFKkPF
GSaeueUZEwvGTGZCnt8qOHGQlm48TD+9Dj14vLGS4YImnPvEKoEhJowS6YL9xjkb9+KVuFwcSvP8
sZ9NJO2abfOGbLGuqN2Pql6EQYgKaIBNwlhkr0FjzzE14Sr4BtJjP0gMO0zRKT7y4w2CZS+Qbb0a
WCWs+hzXK3FPsjdP2ywbaH4sH3QXh6v9mQ7PQ+KJGh4LXdYQPBLGchJgSmWDHIW/IWmF5p7q+xwg
RSFT4mGGvoOPvQ/ov2BCkXZ9+aBjN94Dx4BpPpCem8+yNWxi5BAzoyuloZRMb0ZQ5eNN6qtsN6kp
nhr2NNYX//kPgiN20I5aGqoEIRPeT2lbTcZhOJkE1yJg0ku1u2lKJJ4ul7Q2Rl8PhO3e+E73QaD4
vNSe4lYWDKl4/Egx9TINzPD6iwRDYZy9Tuxvnca623C2/Zir5nr3n/8tMD06bqbVm+ZJakA2AWX8
bQY2MDGDvWN/le3rxxCx2YbjFGjXRqYFEjKmZMW0rJgdG+iuVJDjMJZhQMfi3zMPC1s1OWsmn+Wl
+9d6o4lmr9LelHGbTDO0z5jqBxU9PUNCtssrh7NlONWOBuScrRZ3UEz0zO3OSbPRYMJWO6NRgY7x
jIahZpMYQZbQM8Kb1M8bDjpJ+CGYNGogAx0Cw287Us3WkWkiUAck1uK5BXmPwhtfAZjkL4XuzUaw
xJk8eebdFSI3iEd1wZ4ZKNzRuyznnZkDTLSNB/8xu4H8dBWmyi1C6yaX9Dgj2mBuevoXKOZ33Tew
MFQU2pshG2Iwa/a4FKGyu1d7JH6JaBkdQiMlrlz+pn23Qa8ygm6eIem1EGG6JGeccoec4hAhRAya
In266OYU6UnRCn0tRLioDjqOTgidIvwLnbnZB92fz8ukUykpAHUwtbcrSAiiGxQxdMzDoNEuX8u5
UqETzGXIodf6razcNkG1ngJbRCUP/NheU8pAQVekG2HmKfeCvgUFY6OdovwBeDNZCeIgV1jhXjLs
ItFrk75lX7bnbVysB3/01ET/7EFTSCSQXOjBbIn07eRNy4kThTevXhmr2qVxynDNkr+nRhzhJHku
snCg4dHT6K6d2qbQlKVDUETcEa6ZjHPYOzPGL12yqjp8ccuJ2NEznyxfuUeHpqFfltGqrDBbeU7/
tRC9UBXm1pMdaQU6yx3fMAjwwAgBlROY9xhrwbzClDdGGQYijQaU4wQty+hT8dkwJ4axl5uEEnSM
3+JWUMF0lxd0VRRj5c0rIOIq/MtzxHVzGer8DypVfZh7r+05r1OHUf7jjraQQ8FWUUqrnqZYyjx6
LLj0VtcqNrO6lNjtRDfXMJhgXm7OvE8oDDXsr6seBWaquPlEeAVazCvchsmaIjTuUkHT8+mGU+TF
U2lD8TkgLoP5s/U42JUXvAwl3KLfc5/oU4xn4FYKvGhAEO4DC0yvKSGJB5xWRB4FnhTR4KSk7Cc5
PkkKinQbHUNT2dM39dRcwrIKDlhYnerPXF7Vl58HHRniYnaJx64PtBVMvJe6FaGBk5OMe9ex1mkk
hczvBCWGsq17VW/ARB42PZ7NC91BqhrwQ42P5Jp1QvKstwK1WLRB9fbgxbOVQUVmkabsfVCdpIrU
ghU/4TOXGyMHulEeWijdm/0jNzyQ4OVFK0lPQjmhRV7qrXf71g3AvgdO3omoCvNgu85b7VqTZrP1
QrOw2awEEzzoOMZsE1KL+JlOCv1reUWQq1gh80t9tSPOipS38TbyyBfMMKf7llnFBAAs06adjz7C
5gdCU7c8WZvjJaTofJDliygpz5X8LurSfg4b7z4J3+ISPGNCTdE0GvBNTvbFqZSMLnxcO/GU3ACU
8aVOLvOFgrS/kmeJ+rN+arWjDqgHcXPWRZoM9LRIYbSYrszSyWz/zi5a8MtENfG6I7jJ/RHqyCfi
goUKithydvW0g36YdT+XxR49kGVb0x9saBcbliMY4J5ep/XyRM1Bs1O//i5IdNwTbzjng52bGJHc
2ZC8ilkxhpHFnLQaxjt88BcLA7ulhU3a1uE2Ww4Yvc+34bbyn8KYz3NNCAzCkEfy0KKvYechYZAE
0d2WCKs2UGjfE/4KwvqP6FsR/wjkGIJxvDChTUb/TlB4POYi65+5mupWLpOeSVoXcR6mF0yclabo
oomK0jSSN1OJkDB8RSLKl/ARj/+OgurMW1YON4w22HMVrCo9mm0Q6kPmhFq/W41nG5vLm0NdvYbJ
CNhTclKZQe42GMWhwg0/P6S+SMw+M8ED/3yVCDZq1ULQ4f4Jm7QVBvGA7DyNPyOq+gck/+wJJLWr
B2Ou5+AeZXD/EeWoxqHdnssBL1FJasaPfFEvL+PHSj6FcTUrwmfaKXn7XXvwkY4HapzLg5W8NBeG
DWqHTlokvf1K1uTt+4BW2TuKQeLqPplTESB2204DOpeZ/907zep8k4EKivTWkTOwLDzeW9KENrC4
aCkCOBR97hcZaDrpWqOe8/YkBTjDj38b6cQwfCzX254DGT5IClQAT1N1js8wbO251Quicd+/yXZY
MZSGoLPoTNe5z3C2SWIurkbFX+pMyEnN3DNbcmSHQbF4EjKWbuRnCehJxDxPtJ09DB4J0C9eslQq
KG3WOM2cBRPkFRzW57ZpswYVktq/1sG9QsBZyXwL7f2v0fRKinuENnZT9rH/XcZzpLIAZNF1bP4b
DfHBB34l1uw7Yfzj1uH13SR7io+4zanA3GHekt44cDRR3qKa8JgxwiamlmDdTaTKEOUOO6VFzVyt
PkWk+2a6wiE3yRM7JSt7dqnCdL2IFF8b9k8iECoKGbR2yq/HVu/7G+u8KeGdeE1VJbwjCGh3sGHG
55mI8PbhugPxW+SibhOUjNS7LS45cevUsxuGZ7ljy9OXrYtQYr3vOaF5IrVlEFc/fLgz7Pyd8G5Y
EsDjCRO85w/gpSGtlcpyIxIOUfpO5zBNlvzwbEwZFt0LyHpMaRsuNhKCtQOWknZup9vInz0QuaLm
tPa66RQ5W3wveV6R16St3Vq5hZeAL+gEjYG3OWHPZN8n3RDJ5id+EdCdLeR8LRAig2IbYQn4fZ1M
Nl865DDYW5HVDZDWObkQ7F2cZcCusSorBl0nsTBuZXKPkntxgjzty2Gq8ew8mzs1f8v0YJoNK7hU
OYf3EWuJhKLKP+IFZHzRNkcGvsT7HGJm1VFBJwPC3JosRHQsQIpz6l9rCGmbXUMqLu8HYtu4SYef
mkKGZsgZbFkUYDYrEfigdO/SXTT/UmYycC7vfiiFyanUOHSPdP1I5qzXRAxkrfzW4YlbfpKPbJ2n
chL1Y7Jn4eCNfz9Dp4nnybGWFXl36cz/u+hvzh6AmCy9dCzdhVO5FFEnfc12AGux/WuHQZ91s3dW
wvcFYThDvPEVvRPtc7o5F0VTn3Vs+CjyzSzDcw87JRhjY5gI/NugwoRwfF5+7o4jw8cRnOhDu/QS
QBoE6+DYk8nWwM+vyGDI6nD8S1Yq3weLiixTJ08738XV3T3EFBPPLwQh2RKsaZitbt4sofVcEnS6
6HRx6ZxM4/8eEehZ7/28zbKqauuNpXKqBHbYFAJ6g4zN3eLZdnpEy3PXVYWoR6Hi2hdsXqjSFibK
4gTqg3RpoyBczeUMjxG90702Hivh4CmyFjpw/coN9JU3HIdev5sL9cSkRMZ3ZIKFti4nsXvnWTFA
GOZreOqAAsowvuCS6A0zn7qUeYlwkbCMqtGVMSeICbAczABlGz3MkLTZjwV4MoSZwyozMoeYzIQX
wV1fB3Mb+9bHuIRtjxe+OUe1ZkDT54e8NKExHdBvqbKWizu7Y5nImmlKxuyDiMcZVrcxz2CQaX/k
BpgZwhFusYgVl8ZVeORi/kQfI27SpNUGCUnkK2225OgJdulIS3BHQuuKSd16Lby+3b54ZvHZvMAN
ELJzPlVL4trNwAmXwz8XyqB0kUwhxItM4dLjSk/hqyW++3y8mefCOWMfC5/TBKze4GdTIbzoVSvf
XDfEItZaRLV2tJgUd4VGlGnGHqae3ygbX6Cjy4NB3F4s0YQcxzsF5tKPib0rMbaZjJbWHmUc3qW6
PCZdBFVPP4I+Gww+ORiB4h4hwAsD3OAsB0M6ErmY20h02bogkORkbVzu4XZ5cZHOL9Szl7Fesnef
7BAEjTt4MD6Zyq1gJEr+ZWo97M1RkE9iphJLTRfQv3guZS4CofyJEAFgt5Ynnsz+3dQCK8Tjk2UB
x4KwUJekDKskLICoQyLR33iF1nlILG+FY3vRE/lGH1kCjpWE3KtanajZFD1s36pR7ETLDlDeX3WS
rwTJFiAO3KJ3Y2WIYcWPoT8XgWWJxdzZY2rpdLajfqZwtiQ2kuyao5ER9qJSxXrMSnUTp49gRi4B
ICyPoiYuUXPDCFWv1XOc5K7oCmGp2QTVf/zonzYQd8e0bW+XEwzDG02pz5YtjYZpqO+gOemeCGJ6
AjjAOqe/6R+cMtB55S5uKXch/hQxkdGDFBsCLE8RrEujhZIW37mDZ08O9wGno2Hn7HIeGaAgieMl
BU1tzrB8YIZ94ijrzSphTbS9GVrjcXfq8Ql3s8IHZqZ0GIZRbsXdZO/vs9zlEywDgGNG+KfE3RBp
w8/Q99yyQPcFu/f5inHl40ptyodrh8Dd6kZJCNy/TiAoXMjGZiHveVy6iYO77vOgNBt4ocvR1OE7
JZxIPJqdDmIpaRX7PRmAhH1sNOnaJbdyhgaP3fPFQS48xpknRnXk8BrZpjERQxllhOqesYH30+Os
gS6J5suHdiWwARA2MS7DuNeRTiNzMJ3G38IAYj3uKVeegvT35VFUxVSaQiIea2khw5rHiJRJxdO6
UiswwMUloWas+CpEg9eNuLs8tpxqvmU43BocyW4VlVfCjDXrH5kDzqMdkR6C5/U95FMZKMudmp7q
yxKPoK9DCfdrp+V9lixAJ8v2Apu7gUA3kwlDL8dddCTxZuhe5tdRl1WQ4jplU1A5EzUHavaumo/C
tXubQND9WvL5gbrnlZUEB+KxPg7hE/LoonQ0U6R924D8ahuqpTI2JY4NhlPVprjDhMJErdv/AfMo
/Doz9xJP1m2LDOr3MJJqvcRhB02P4M3MM77LfJqurr5z8EDEAICFdM26WzuqpXZH2pRp0ANnq3lp
HMVCRlT62k1eu58LWZ27cUE4OBhjLF8O8QuL87srKioUVqzKJISiODFS04liygHqGlAQBzSp6FWQ
0LOW4L0/jZx/widaRvmXvIuB30rXrrEojIMbl1CteXrYFIQdY7K8kp+iTX9CZ9rOuEr6j3PFG0uT
NfxF03eJZw7R3n56HHIDXvXmVnLCyZrryocDUFh93aM76phkLQeXPwiaRqPv0tfFlCS9OidPxAFx
I+nZNCObmzyYjsTKjcoRZEbewvdSdDo4BPo8qg033L71T4Rr+5FOIZj9MoMmEIYBjTngyvd4SK1r
FrWU/UCbCiS76MQBR1q0zNsf/FxUb/STd+yNcn37PJ7ajt8lsG55zZA66K/EHNqt9PpmSt+vCO/m
PovCEnvZG8ZqLNdFc7S/3F0ggNq5mUDXeMUE+s5UNwDdXLNr1XM1rufsSbsj77dFEEi4X7AesTfc
igkRP3kAfghRIUAD6u/L9vps+MRO7JeJhPw29KFL1VqikQ0YGZ9WVyzJ8IFdaBL5imro0l8A+DOx
heV0DeMYxuAhIXwfINBH7X87DokDSVhPBA8U0EbB9WHFAnX+1G8vLE8xTE6Fo3WuwSwibl4rRmyR
7nuSNgZSRqpBifGtR2OueH/Wtyyu7MGlg2FvxQBB2SojGmGfcztHVMLUEJP/YhdNbtB3MP8kABv5
VOjqByEe7yM9+VFbVJC6Y15dSxqZK1HDDlWSAZj3kX27QN2LfC75mGix1KUcrgsLpzokECPwesVI
UynuzAhoHnEyrUPtZSJDav6tiWzvirDaXyo81WUSsm3VJb3M36DrZ1F+cF1y+l1oCmuZjBTzVboV
QAJV7R2Kz/NiB+gIvRNyPDd0Jyn7X4KFOTcVbjM1QX3rW0B7gu0v3xwkfKQMKvgKHl33omawwW5V
EeIJpusR8q5UagZ2jjb5GwTyQpJPaIqP68QwlkeaOyTjvEQ9Bu5cPY1iShMOCC55F5WxXWuQxfPU
7GtPoD1HyEAvdClFFvfnnWlZunX4F7zK/jKe/xUJq2M0Aox+UiYHOkAnfilLoBhO1MK0ZgCwLzsA
XIZXjrCUd7yo1+JIEtfNEeJ9uRV2va0ok5AlxoAQ0eTH2GneoFKPEEebJqq0m+iXZGSsR9i6bPOS
SjJBwLBTBhBB6JBbS2TISZz2eHYN+I2KIiyi5dqDiDO8V0wVDNQR2+rZu2OQM/WSRbMM7uGlNjuO
KK60HXTfXum6adcQ4E4a2RO6dl3duJwJssV/raFd5VjZqR6FytdKNTjxYDHwbndIizgOoRENfHCT
FULkI1FDYweq5aAiTfPEfDO+H3B84p62KS6wfYzGukUK3NhtcLg3avPQ5qWo/m6glAFnB2rs2DjZ
fGY+tFzvF0seDzsU2AAXMbMwpgjx0WzK8MqAhPxZHYpKz0cY2W1REt//ILcpMd7eY6mfTGDwSdqB
wnjKMS2QOvMyrF2WxgAvKgfm4OP7GzNltC/vPMgNHn5quYFMXQFSY0AE4hMY+MmBFAxnod2kEHZj
D9irEaMhBQWY0R4KZdsjFfD0d26yey0J0g/gpLtKgU3nPBWshtus5mIaAw74fEzVPQEaEaJyD/rm
hMqxtI5hbMptXI27euKHw4QNwIBe8cxgowAia6WS3QyOcxT56giFtMY6XQz6nbTv1GazwU6h/PRK
55hqdaM0G3eN+fM53naRHPQgl1vPYvTGkRC8naDuXscDNpeRfYsVnB3Xulp2CK5kTGU06gtBZ2tx
DezQVTkAV2/+iBzM5X6DyIJjg83bzdN8zk61EBfxkBlwoWD/FxuAZ6b1uaxL5LkJQrqY0pLQsktZ
JSd9vHob1VlOF41snUlwEkoCcqiDIgKMAfRoYTmj2QElD7j0uw7rNllvytCQFhZ3FOkcaT5vcK8H
O3Rh+8GzYh36cq7AbI0M2nxdLZJ+0AwpqC3/LMMDoBNkTuTEJnh/c6Q3WUekVfCGZOHOZaj8wqeI
BokoEU9yBxqaMAD6or5BDkFhoRblJxRxPEzLxCvCgSQNvIoPeImyJzl05V1Y/gH3WKQfER3GvQbp
K6n6x0p4bfwImJAJ93BSVqXi7v+RXBzzjTYjJ+5dHebQleIDLBEudcAmEmW5cKFjO+dzfj1ab36n
yCXh7aEk62LrupfI3eUnx6Xr+OkbyoP7547RwW6/nwy57IN2PCNTwMqkiL6mQiPhEwA1v9XZzSKX
RoJofZ69JgUWQlVJa+QcMi+5H4GI4ga223YlBFZ5JVAqlfcA3CZhjaqlB/7wTwfFMIzFLsxKBpp2
+Tm/0qf9LcmkWkrVIhN8Vs9LcL+/B5M5b8JcZ2kpUWwiy2G/fPPk1qtM5ienyd1vIrvysAb1pCNR
3L290RaK+7Ue0PlzJ8uYB5FFv5I8+FMywh6lbEkJmhXL4HN8+LbAcNbDh9OMDqSePWHGcQ6SHfD6
hdrYTt8HXB1CbQ5fQWtZfBMeQee70ipgNi3DGMvv/BgrI5HCEVWBLmtne7nvjtVjbc5thlkPrL5z
tncQlVAIo8rhGJQ24ZWSHX9frJztv8F+aIocLVCZNLkAiB5mPGVopQ3AMAH3MfLBbnw8CSJhvCBU
0DgKJQfUDxBGwYbSFmnM/k539KDv0hyTl843vxmJvaim81h7xnzfnEwjJK9x7WHE+vf7X/pCA9yW
sa5nLNnJVvrdXpYXFUTNns+l87XM4vNiTXjyNvQ7AXPlQ87YxWEYrl8GMnJkfEFVWauWQ33Ru/E3
EVj9wBHAH55Qd8J34wsNDmo7eUiB5BQNPpCXdhzGgWTPMDoAljWyrB1vkmFivpGM1amrhkWG0QM2
bF2wbco4BhM2GJkwS7kxRETDLZYHvc9vtYY0xOmhC/q0zQizPpts4lDhfOunIHoXq2n3Q5GeNU7O
R3uvOyEgabkCKWqZiU+VUzQXJx9Q0BfwbfRKdFZnnXuaDV6Jl2vojN4rFs2lJWUXNWX8wwK7QyM+
195Vdm5gwZ9ziw03iJ0p6Z2YFjk9xqimCu3UR/NAoP1uZqG4Rx84GyS58QbqNRpyErVXpmnYXVsF
Ugj9GAPE6Z1ZSF0kAo/qWYGkYxB4fjcSxwNrbhBpeuGEmTC+0Rdmj7D0/eOsWjXptjAtH3TJ1DQW
1QKw5D6HFNVjnvyyW1wDjtsOMlj9m+pPcCjnghgdq87Zk7EvA3I7KrzR/CetFlwR1Q7PCWZAFs8b
x+P997I2dYX5212vbqGY3+kYBWgKPBME9P35Ur3vdw8CCSKt30p5M2A+bx3Vu8s3Qay50AjAWl9o
VpOfXgeMDJF+EEg1uZfG4rfVNsv2veNKOGDb8fgoaAkowwLCHD+icc2Omew4vWiUaY4+0Da4lCRx
86mB4YXIyuHP6KD4UbJ2UI4Ra4EVYoLRIZplHBRIet2daeSR3GlKVxjDwf2JsdRSLvfvpDFoUmW4
M2/HtmJlElOrMigVRjdxTWIZq8Tj0K+q4n3crFozo48AJoccjsXmQbbZcOeaUYaF06nBPn9oekzZ
UtIwEDoGwmUdYD4iW/uEz0+vr3D3vTr5+mx8+xL6R0NV1wf5dAZUswy1QY1yr/WYR4bD4SxSCOa3
U1MZCMrtGlJAvFy9o2r6Xeb+Yf4eMnupM9ugoeUpgamLvlbeOvrQn+XHYVIceAmGGTGIvcgRuF2Y
/KOjL0TtqFkxsI+fBHS6mJTEqcsgelVKCqYdjMYj8/f07vHwC/DbC32zeorQUIKE1fBtIvK5mFQD
8qKJRDQfKYpJDGvZILDckI18/d7I2QpbQATBl8feSrGV8BA9WHuuscVGyvlJSMiKtNfnvPr0K+zs
7DW/PgVioOxubmG2620oeHln2JDAM4IVVsLOU4yeC44KIu7ElVmOvqm1UbRBSGIXCXiDwgLjpF4H
gR/onBLP+YRzeFGdfHwsu0ZgZdIslBcrIS3bGjjRTeRV1tCf0AqDJn1GSeaCm64j2xmVXDtg/Vqx
5RkBiwt8GcA4p19VQcpsaqeNsvEGfD4/n4ILgYbVIjeBGcn4/BsIGx7hA4NEkrFqFCGtpkzIrHyj
fXcT0hh30KA5CxshLeXKvRmdFnpxq2vi5X2REU/2V4kekucVeRxE0ISQ31d858YuoR3nO4p9nYC3
XDI27jymE9py4BuEkhisjH9AB5INa2yVyCPYLXnF2mvusCFTO8P3FhZPuP6jbL0sDRVJmPo8FeU2
MKEKw6NA3FUXgCYTGYFURrvphlx5hqMjNGbUd1W3FiP78B2yiJ2KGDS6ZhLsUl3PK5zUeAHbn4sg
wGlvUo9zO+9yZrxGmYp+oUVzTtcQkamCLBYcpJ594RCB1ZMCjTJtWy2GTEeagTLBoXJyautGLahR
4VKhWFRapejt9MWLzSgqRwBMqxhYZynzWsQkW/Kn/eNEvlg5GjkOeiXV8M11tKAR1638eFppxZPn
Rqup0n6/0kMyjjWwCBr3uPY07nQg5WUf+fHiDLOVnyjGugXNN56iFr2P9aygTmjcyqT0kxpDz1A5
G8FovMhE0YMWyRvsRMcif94vr581KpORpa3ddAwAfb28RP62/b+9TRStrd5BVC9UzVOizEj85Iub
z9NbE2IiS/UM3FsfuYkfrS23QXJFfirNXMm/vvreLANrBrC+85OukODeb/qX42XhXdw2vh4BTso8
ow2f5AIk7lnQxyj4deOqm5ChoG4f9xu1cpASPItX35x1M6ZBjp/QDe8d/ppQjLS9kWyaLBioce3J
6nfrEQ5lFfoOH40oBsU5Mi6VsKNE0LDcyFvaehqyTm4CRNVc3caCQ/i5Bk21OGlI2wYUGmEC8fck
ySqINxt3IMfjZq/h2Aa3TO3R66G4lNjMnV2AwFFVGHDDj5UhVfPUFcOGt3GPU2JzcB7T6lde6U9T
dPz9579Tz0q8eFrTH4RhcAMfOzUddNAn3qNn+RGcOeiDDxhhoO3wHo+TQjmC7nV66TzF6Frz4Hpq
uvs0+VWsiPFCag8Sajrep499Pah0HM9WjWPy8KXVKfTjSa9LwFrNmdn8ib33jvX4kn4CdofnrKBl
4YjLFQiKfc6RrC02Hr95rK7yKlWjLQj7G+owKeWMYR6dawINoMLg0FG+my+9fobgoTMmGR1YJPTu
q7wDFOBQIZjXMZ05+inLx9A0SCCnV1mZ2EpnygBlU9eGWCtdFpvAcp6cOGbUm43LJfAwX2F1ucsT
Io5ZeSATLpyHh6v+SV0vQ9bnctV9d2bq1sdtv18wfgi0IXOU1YNgen6h2YpROTMDjvGztTteb9ju
c2ux989nYKiIPstBmdKFlLebAkgDdq6jh8Usk2gNlZW4DVJ+f6S9wKmyeTbMp7P3S8dvWYIeBZC0
ymlEFdDwXVtlimeRbGl1licNAPfKsUPjoc2E0L9Rt6fX4z3OIxwkpKOF2S+TItR3+DfqYtZpzC4g
m1bMwAjFl5kla3HAQyHO7n0+a0ttFx6o6d0jPPURNiz33ucdXHIXxLu1k1nT8M0Hp9lzj+bqX+hs
cpuu4Cz74BRTR6i+xPZg6vXNu2nhs2Uuv8sKN5GMMLGtb/VkZeLWcNtiOcy+ySU5RZAlhv4WysF4
DBaj/5zVu0Vc2jZpX9feKtC7jpkBjhgJnC+YVM/hgYyWSLnMGrZF+pGkzIe+q83p1fyjSudrW9O/
6Tmsg5z7xDCDh4dh4v3qrrMJLq3ltr4V4cCgiAV7BNDsw+F+IZkOxZsJoHppvgwUDqoHeDlLAsDm
W1kV1LS18Eg5FaomrcwxUdU29nZK0MQVQClycj8itXfSoVsFsoHAAVCamhiRgctJX7z+fbMbXSdq
nOkR0Bm8PrKbCz5ZQGCKOvOZW8dF2LxD8xsOi+t4qOR+e1I8i29OxEAj+iNeUhFRuKcDssDPFN7d
BcdAqfOu5oyNkT7NURDqjW8O2/pZGJZHO0XeqWc5nReFFvuGWl0VUrqEjA+mw54jUs8rt7fE6tnb
ZWne1eS59ZFYZkfuxSwCAnbI22qxnVtWspqBFNvvXE00B63y9VX9HKINHnn7rnxMF3MG67vMfmW7
NiPc+pqj0K2ybZcSGreZavCXFA1TtZsM8rIqI76l7pan2BEDfOKnMhfCkdPrRk1eakZ4BHKXJa7M
2GAcZ2euvOyiKyNV+Qdh8/omg5l3UHbCuO8xGizYLd4MfzC8uGVzTLrTFGXap18+zfm3du8hjgIr
ZgMam0UaYvPpwzuJNFgE5b2TUjBhXODajApdRdXSMUp4CtsTyD5StkYYjGDBEpeNol9n4jX+Wi8c
0OvkN+8nIsvkaQjwUx71bA9gdaMV4hoQ3lazAAhvSOmmbBQpkNd4CC8myPqaxIW4d8lccTyhxmNo
SoC+JbME8VFaCEmc6mRvEFhj9Y3shJkJstYWf0vY4oVHkB43RsHB/6abYPcBOHiorbNT6DOlqond
89FdrWYa9Zt1HNiKTQKs3VzVxEfchHZhg2vizV/3OndPffvHBKgeZK6/Lf3qOHpKLR3AuFDGDL1z
si1ocdAWlxTuDLsobGUbJIO+XDFzO1RzHLvUPGpfsFrKxzzc1+UmLD6JuFr82zvhAj1ij8OrADf/
IL+kqtRuYOH92ur337jxIskRgDY6qKaD76ckrj2txo7au6poJa2k7gCeRFdN36UB6nwSXF+UCGVD
jcoavdP+STIbc98aZIev99sPhG5+3nxf6kd+RI3uEeaudBrDL1QXcuTaETCBZlFW+vAB7/JK8XCD
NNrfIeyq9V3WxhRXdKyLQkcgqrLE5Bn4/Jau9915gPdFeKeoLBwBXFQyiie7pxyWgPinwhGRM01a
T3jVtqUpTk0KjsP9lMTtTyZPhfc23LehZeTkSbcqvv36pzYq+0CMu9l5Vch3J4nqPpp8JH3fxvS+
wJPqJBiRYjiVWDbI3jJBEue5la3mT8YVUrghsNaUyOowlNW7AmJ+rLs2L1ZK0+f9dlan42BQwfjK
dI7w1I5ggrAS0iyq9GNgVDOdnKLUAwd70fGnIxFMoCqy5zwmXaA+ytO5/G1XpEbHoAoOxMtsHyDk
m/F6uFgUzM/fUCFwFOu4HTopYuNAA2t1US+JmZ1TzRAkkZszAXUL5YzcUmgDwceUNJmXZqTeC4O9
RNP7i+gQSi0/n+8PrJoN+6V7NnjYoKfQx0OFH/eRCyjaQrLURLSrKSYU1O4ZWGmH+U+UXS22re9h
4OM5r5D+4Sd5oUD1pdDis00oMTQ0Is0gseD5uchu3CALaV7q3ZxJ13KXpjw5TReJzHFGhY6atzIt
XjsL87pbJJo5CFqwWxM+YEiXhOCVtf8NKDm+OIu+u6Q6OyLGtamHYOBGIcMZlNkBQ77CV0wUsRuD
ub7bts6bEGWpPditl5iUV4EWM+8clKNnCe8BeAGyCEmg2MJCQfbzbvRg6BQmbO1jTMb4vCkfTpxS
ciar2XTEhCdvwwx4UQeoOiRTtA7xGe5rzRYRTm6keLxfw16nZ9Eh4Cew+eC3iLXmncJ45i58UXvP
HP8g/Z0P/7kCeKrJ5q073k5NrERG+QiTrqjNH1kZYaZNpeC0uN3+qBg3bCwWBGIBssEFf6C2/zB/
Cl5Rlu1gxhmCGn80flT5OBF4RC/N+aGF5ag1p4WSfj+R17kWcB1FeuSz0l2UYw/6bSgSuCpcTyS2
gXFnKL/8M3Stn7EvS8LOSmZ7Fnjpa45lTUqzFHSPKBrXFrSQ5gsTVuVMd4RJpSMj9P7gp2gTHCeh
4JJRquB8bpHgv87VGJwchUsSMfTd4XNR8tLmMSRNMjoAD8sITpc+hnxY+wBZvF/MBCEzerbmCDTD
/mrP9lpgt+eGQaiugNd3UPRXIZn0VVKB8U1uCmtyI1EWiTS8gkJtE7Ji1IXN0BwpoVpMmnDornSz
zsxpJsfXM9RqoZa9+BtDxPRtGx6qqpOZNYe/K6lrUxzLZ/KQTbxAX/AXfbt7QsmyC5A65iIVtDYP
uFBvkJ25mgiz1wxbQ93Vuuw1W46cS14tULduhWxUekpTJ50D915ON2ic7478vKwgYlCxtcwAcKla
F/AUPcRCy4QclrsNSF6fU6yvCbqL4Gws/M4msPMnOUhpRFj/yKmCMBpqyIXABoygdaGBBTU5Ktoi
m+CFMMaivJWBRKThI7U9yP5yS638djyRI+bQV/31Itwnips0FB9tdy1IflscBLxvWgazneN3a6AF
sfJCZi1HlFyORLp1WaAoPMJyJ60w0cZNzERKW3pnyPf0f6mCY6uFEhpM16iC5ROOEaFLHuYK/j5J
hpELqA6al8TwgC/H6SNxW23vaR1XR2MyLFOvW1Mc0GIqX3WbQVzco5mcdQBGSbOu5e+M0AmyP6cF
U5ky89RDrOHpVnGS86ORU1vDwHvlLIgQ3ip4nEjo5tbOvYLxFo6goB9R0/qorD4ERPcJIq5R9Ckg
Z0ar5/IWDdY7WCnJvAoTi8lJkr53JUmwvxUenLb386qmTeNmjVTSMrOgGnqcHZE/mmbBiBMoQjgd
q/hjPF3edRDqJxeaBPnVaN7ahwU02gMfpJm7PNIWjAJW7rvud/zpt4v7CwJsWDoE+8iIB3uq1ZEc
h5+Jvvhd5xfWxDm7PdhO5QV2QoaqxYQGNyEelzkVzVHm7CM3Zi/JSQ/MGYtid/Eme6iaOhxeJ9bz
VqMv4C7Br/oFYtT4NWzAjPH/j9ah3i+TlSXAXZ5zYOJS3eAib1TbbTh9sK0rNzsBDnjMQWjmdKmP
+jzGQHiOhEw+tw2YezUcK7iWHrW+mPe8z/i7x6vpzxHm1LRNmkhweaUJv86lAGmVMeAOesKlxCEd
1HtVFtqaXoPss1jc181T44sJfhSaiqyvIrOThx7QkT8KXqKKkGX4C8muLdbuadGu3ElujAxZyb4Y
Sbb8hDiIfdNj1by5D/eepaBp9jGo1bGicomqjmazEOL4cisg0ESvb+w7Y7FOdZnZu3Z8rW8ky0Jh
A4WA6LbZv0tYgWFDsBssvkTGuzLck6LBS0ZgY++jl5buDQ+XsDeVmWUUN9m5CdEUX6ZqXqIAfHG/
5n4q/F/ljNM7yowodoX6XyEaUbw7o6XRacK9EQsEbAARE8StUymHJgztfidhWn+N0GGMLw7/hBj/
2Hv6BYZVruE75V79TF+xybBYrctwqLFSY5BirGDY9Nfxl0R5LHfKtc2NYLepdCc3SNKzQQeA5mmD
t2pW5XCZba53ywmV+IgWr41BISl4jlUaL60E52prLRXRC1KsFsBG5a5yO4H/UplF18lCBPBaCEWT
pK9OiQrdElHYWIBSSyj0K3C64Ux7EkuxV8dn3RLzJrvdunnZnY/TpKkn3DoFAT1qjavWrHoD21pw
pEtcgGIXxlG0CUJY2SkO0bu7Yke2vlOBsdqR7RjDNoL5L0uZ2G+aN6mheFBGRd2bVxs3xTnY5bPY
vXV6aHUe0XchTizSjupWl+JdJI8aFtQxGz+SwlZO6INuf5DGD6mnhLKFuHR8ntza45sDR90VcrRg
BY856Z1x7fivKHTpsAf4PHsI4emu144UUiLOJlBXKE0HAWTO0EwU1QNPVpyIUzKBET/M6mGd2aPE
ruSwezxr0eXcyMre6e4KT+Fn0ZwhmHaLDx10VZ1FWc0fS77iDpxp4nLIYumwZPagxw3iKJRIcf3+
UXkt4zmxif+QOuSFCghXW+P2mTRZ12enDVgra9W8RuGJ0J1QoZ+UKVnDCFth5jFDPscTCMldZCeV
1qCuCgSy89/H2PAAeImZqeNWPVYyvFeW4jOJItvY6Xmr4qGn6zlCPmiRTsI2UrUyGTzwmVpvDJRi
wtwcLXFUn+RnTQh6wAAgTXrS9C5sLwnTECHJ95kiEijbpf/qh3YFtXp89sEdMn47powo/wZt2d06
lrtvSX7Xqr3GjvUcyoVGIwc8TiqJK9AqR1KgnwIqeIStr4bZmKKkYkSjoFMN9Vxr3zHkkd7r2p6S
NJcy9J3X4Lx7mjxqXDv3wktbl0A1ohw5daawQAAnJRKpZp+z5qytqkq/Pp80h/hOfJKDwNw3h43W
iE7c/0C7Hn/vYuhiF7MiW+p9J194GgzRtVGW7TZ7CemjLo/pg2qQQtsuhqi9hIYVtZD7AVRURH8V
euOvgkV3rMfi2iksg/so1ZkvfeX/YWRekTR1aDweSSHDb2XHXF0gEa2rX4QawnTiAI8R2gHbiyAu
RRf56n/WrJiOAnCT/LosniPnpT9Vo4u6/ZCD8XW6hL4iNbHk4TMaeEWArNAQfaVwyM7J2JVvLXW+
0zxAAOZc5o+e+bmGQvhy5ixX3UaiKtnNMIdJMPn1AtY4v5mhSE2ziM79ltLtjKKICcghmft/AuBN
6ooKm1x+1oTip7IXqypb+1DeBLd9cR1my8uYXsnp0P2Xu4l3HcjEXsOQuxUQ4+hY/9wdBYr3UbA5
syvuoGHpQe2UlO1JeRg0OT/312SqyyXFOB+Nqh6GJTjkJPanW8EhEsi5eqPEowls/biHUxHPlp/r
VRRwp6dLDmviHJQwgKIBQ4YarctNdduq90UqKWLM+t71aVxAhGOhiBrmMsFgACYweaff7gwZp16R
neffiq4Q2OwKnE8CEDhXq2a8BtoAPbkfBTBglRqdzAA1b6XNqfR6voLZqYQQXSVBv4XeWrP0hLNV
aIElYqjn/SfYME74lbE98t11sMloImVrMNkM7vUyMm/XOs4NLQTigsfK6v7/d/JaEEPq2djTUuvj
1OG2cj61dej6Zm5ZFVyo1Z6GeCoNidNaiM/6tEM30f8wqYLsXD4AdYdBbUwkg4qWOWtkKKrUaXGH
TS2J2EElP7lVXrbRNkCNc28cLQrJ5FBzYvWyJ2YSK5Y/NMTti9RA59fLYrubkP4oy+hgjE2nLaPq
qISVNWI5u+DQFSJGpuwAB3GqUj/dYRhUCf+2sWyQdv1fHEgGcwQU+uxlmqEEI3AlAb8ZUw/sdToy
LZ9PDF2uyhKqe5p1iZHkF0Owsw4JWtHyL+nGG5moC7aG5bsLfSbZLPFAPMSyzgulPKU8FMrHILWA
yRBEaHpCbYfmsZ0YGxqqRQhtKB257j4HyAaUzc7O5b3PH6y6bWaJ8Ckh2YohU8qUDGBgSx5HgDt5
uR6LqKv6h7goS+Heh+2YVAio6pSTFk6v4jocnYH3kDv58vjStG+LDRCXTGE0YJMvkqeD5mbskg1P
bVyW1nRb7MxIzkqkezd0c9lgUrDHPrvEuz98kM1+0KGNuFpIbnqnbo/kT73WOkJYm6IfN65a8l3I
5zDwgHvSzVXZxCLGVsP5y53Az0TjZ/sLoTO4NmJ2T2RmIlyPcOEWBkmnu3OJ3XRy/k6S9qTCd1eH
/UbEKIdgeB12tgWjiQdC3bFWG58IE450Df+jb4XZ6/Hz1xAcRTTGGFUs0Fh4dxQ/W5zt1gbO3Vrr
VNHUVu8dfo/cA7UF+by9gfYuzqirUP05DBboJyE2uJHTb5qQZoW6VzHPLYrMgOKBqjK9jO/FdYhR
sdyz1KVg3utBSg9vrqTfuDBi7Sg0IYtLrMCS+nsQUE3LGPgZGyv/hmYI86ZeleMzO+JpzLiGIks0
6qkj8kMeOYX2oEvwzGyNGoyRcVTdqlOLZbH3GQUi1v17tBsfB8E+YjkX4mTVMdGyacqT8bwAejOH
ma/O19fupoixcC+24X+BX70hIhWKKzjm6IkUA/txG3KfNOKUxQ/O+3SJ2UGGboA8UbCFN57w6bKK
Y4czlBj6d9ML8z2rkjTCD4ZVXNMWVr5MdTti8WuN+SJkfc5PDp9anV7qOy5ga23WaGGq+ptvopwO
Q51ZMLh+MFx+Ur5jKgyTw8tln/rTvP9HOkuGDe3iKK6ugyGizUNO+1sbV/CFJfQqGffv/xiWjUae
T/NFEnxXQm4ILcy85e5rbjoZ3VNHbLvfV8O5ke4J0veKODXRVsIKynEs+TbQF+7i9TJGIcfj4p5P
eGf8oY0gcvdhfWvvohYCuwnB/UT3W+gtXRifpr8TOqRxSfxYx7rHX015txt+rH3YpyEalH2+a1Me
bdDsd0HYBgrCtgrhtcQ5imBpCT6q7GnZ2KP0TiOG0fP9GBBD4Vb0dJR+WYZBbucYHaQURPQxGGfN
PrrFIYpBiphscvFan/fdyzD2mHDBJ6+MbWWQPp2fFcSRSeCbnbAom81dg2piicEGHhP4lVI4gsY9
PHntkZ9TrQdC3JAsW/5h8DJhLY4MTkweZgfBe98cvwumLGdABGkrwh7xmVnrhTgZWUTjdQVMkqxO
Cod4VV2CVxNaDxvMbLuunAS2V4A0dZV1qS7o5LVEvbHeP479TKL+cF7p84nwpmgBj/LN5oIMtNSm
lNvWod6fTHz2LxDiiIl0uwMrFfQnd0wRtbIAME9E5C7jcnV4VjWSzbdpGMY6llOF58WTBaPxyB+R
/RCHpzrRMgH61mUdCAehfYt8vH47cEetWxneisLsqqKvG72Qm3sgYMlHDb81qyAnPWuVw1T3iOZa
AvX+u6qxOXTihuTqUvc9seJ67imwa6zOltUlglgQYWqpPCwErVUarM8s7GYKDSSZLc5sk/suwkSY
3NP/mTnr85i8lNwBO7GeY6Ly1KXIUsoZm9vi7+4CL7AONOIp7yXVVBWBVgDfN8EiIU+W5PpBIxj0
lM5ktFqMI9oJ2yV36NmF8NrIo1k51zykVwVn/licXpxRXP24/LgnGKSH44P47qCci/6tZfm0kXeP
3vH7vpa9lZAbD+LAoMtEcNm86OlHm2uJDqvUfVL3r6XuhOfDF9PEVS61YD5bAYp2akFNq9thLgpz
sBPfpHAipOEafXA7PcWAL7Pvm9cQCl5FZvsxqwqiDKdPcWK8QDleDXnm6VjJZRig/byoOUhcmrZH
qr0eS4bxatbI2QDIzgLEZQbYH5AoPDU9buwRpN8YFi5C5PAPPxhoFL7cS/fhog/Fvt5tHIUIWT1X
w2RlnTHB/aqUe0np64O0oMpDSJMQLgCEaRXKn91R7EbxpWu2J5a6aEQDND31Koupmfey/SyAmMuk
KdoHUN7/hn3eb9ixxzxl+ztBD26nNG9qRkP8Eq6cJ9RTdmGv4KXQejw/g0naz5vARasuSyCR7w8J
MG1PpVJB1ayBzaAgdj3G3R9KGLrhFz+/9aI/r0i6sPAXH89d6Nc19jheRM+BA78sYWy/7oCvgbBN
QZqXNn7E3MGiFMA6zqUaAL/BNxyfP79KnSNjyevKZP7PntgN44g1zro9iZRpcwzrf/6DXEP9IfV4
kiJse8jtmCoWt4mep8qN8cjWOpn1Qp6NaXj3yenVPU4cR6I5heu4Ql4nHzsceZ1ir0rFb8Fi806c
F5aKbFMjL8N0mNDpuSy1pIaD2VmfPL9vVo7bK/GkXHPdClq/DZQ8JftYUeH/2A+DZr7Csy/rFlJm
0Ya4V0JT3cboxK10whrrseBZY/UeoxoKJ5yiGxTLNu8TTr0FVzGXC+6qlBqTjcQDgz74VRDKpFgo
C39wmAUMWHw4WeAPT9iXGW51+0FlQoD4c/q+UU3LDSs3UwvT39MdoL2A9G+WFeJ1PuOEVNgMnKFD
rHojDsh506W3S+cKUK9UrFMbYNR2ZPuHlCecilwYqe+/MLs/45+21EM8balkuYRwUg+FpFwthwmV
l49cFIY64bSfRi5Kg+kor60L5MB8mdRZaP+oWhpUk0UD3pKgdYCIWucHKHLVKYdeupA7hmJ09C7R
OIblGm0/wztPsY+odHIVMNFmHlHYiyPLPbeAGpPgw0oV0hGbBMHk4uWUCuJtxk40TQo/ZACo1d9c
R0IwBy0ly4ganHN9mNCkVtlizhuqB6KsBA32UocPgKWlrgnlDKhpogpbedBupyFkvf+HhWLboSuT
lfbhZH9SdnUtJVR4zPCR/vib/1+HqVC8UnSGkRviiN+RsvLwhAERmdRWl6aAs+kpgEm8ZgYYcyTY
2uzl2pew/rR4R88y3hYfe99gWqnh+jAKQ+HwoI1USGV4gsDKKnvpfQmdiPoM0DCbYsAHZIw+DXX+
TFdjuaoxlGKfSxARfn9IvuCUh5c+KRlMDtAQB0OR9ylxYbWAzmkBttFlohLb9CUeNtX9yS79P7cc
dLHs+kUQt2Ukve+I1nTB4hKTyDkv50WpTENm9V06ku/983QOcHSrrrr5TsJuDn+NOLRjILVqlizw
XC0xIyHqTwwow2OroQQsOnt0A3iXRFPGLVNQQnRReFXLMhIwkQ8vEy50RLaI6TYLobmP/fnILX+b
CUncLrhi5HA/H/mJAtjpLD5jdp7IdztZw/b27qdfdgpNIbsUCwR32X0ZSIxwgtwp+ZqboMkcGeJM
gbfflj9Ts+cqKlRePGBf0LLOytbSy+emcGiwrMWc7ZSOAmCERCJVXYAamBIjdSxGaAet2lXC4VSJ
J1/TTqQSVx7DuROg6pMYLFMyIN8e78kVyMbNAIs6ZEjPbdlg+ox1GSYjK8pwvBOUJHD8dT1Ti7Cl
uuXrwyLG2pyJd4QUinzD0JG1rbDbHNk8bv6IbZ23zztra7q/7bJyf9sce0EEcGruOJhOrouAicHs
EezA4dgLmZjq/YR+JRim6DPlWMRVLmLbF60Oo2JzPQO5VMF3bm6wmUhN5cwVBUqJLppoQq/Yh2b9
zSJYF8o+oYKSJfgQN/1gjLmnnLWPTj/P16UYigctwtzThmGRRZSRALxm2VvLkl87zaMsipZ8lHFu
8uaNlFfnDv8/nZCWNuMSzi24gKMElj40QMLSU6FjsWLXenyh4Q/N6BZjzrQwZ8fhlxRC8/RvBM8v
Q71E1YAwDsK1M7WpmCD+LOzrsP1pAF2m9lob/aZb93110PXHVcxLoBzUICLYIiPHpaqaiVdlbaJf
vyUSZR5dPehvPrR//8EqtRdcU+srH52eHFkBlv4lmCyNuyo4DhmRVuGFLjNWkAJlpKpwvKVDOx4/
STNzn5JFbMejhbsnBsQFuGBeC7qa/WOQvjrIWCLv67lgOx/YPeD0KFyJYXajxTwkXFUiwkn5258+
6D/Sf6qUNXqWemQbNa4ZVhrpkCXYfnrPblsuERHUt8+YpjNd5emRQtgBtaD/tS8fi73amhpxuc6R
w2r/YPSzAaieXmrEaDGRqZY3JMcCcrHzQIZATQi8ARfcLGul2Rw/Q8qlkQgqTlYQ+vrR8wRZD1fZ
bq5/SU/rEU7NFBJ3myCcsajpDhwE7EJSyu2moQPaIsjG/Vwp+QbitWtXqe58mpVoWfOLLlnIoCBA
rD+cTwbQVsk3kTZfqUG3GVaNmGMjxkvUvNRD49iUFxQV/uaRFzykOERi5GgDLikz80rEf6UcbR31
EfoZam8Su58rHY/DvXjvPPQdL+cIV4Lu05+Bi13QWLamd9rdTSz+XDTB24bz2ADRdGfB/dW6/c9/
lwTbOX5YRsx43YAR3YWLXbyq+UYPB+ez7uikSlOfRM58qlVM6u16XigdP+GSOSmsJEghVSaQof6q
YEz0aaya1rL71prkvQZohv6mbYO+PGH7yFE+MgB5p9cj6Rw21yRhTWzhUNCwlvEto7v2dThTRZBp
+Gr4ZvhuejEHYsGGrBNuYLj+OXZ2+yggqLyC6wS9io7HNkiXof0A58EjomRuC+xY0lyQzqVfpBWk
GszpzW5fY597bBa3guUnjDhJmBDSlM3hLnXBpCiB2aP7NAJvFFsOasPUulNKyXM1qiSfRX1+bdnB
tQWiGsvBtwdz+S+HxRdFH2QD0cUCasWkzRpEKblKU9Pae39oEfNWqRcV93NFvM4ZZnlIRIjV6pfD
HcgUM161fL/Dzi4hXehRwstHQqNkEv9GAYpJmBkM0BjyyWB3cYzBfjANZ0TeNHrFJ1m5+S/9O92T
7AbOiqNO0ZQxaNknkXj3WsMhjHx/4qE7CZVac6tFof5HRnFQuU6xLk5snNHDSLPTQCW0uzO1Lc8x
0GI3tItGiKgnHVGaj+UaBNp/94+xB0WKVPsSXRVF7a2OgEdMbnGr1n43hp9d1Ezrg+2RfxWtwdEy
HcLT8EXi5lBTiyoChubAdE/LXjItGntXcfJ6CsWFTFVQGPcq1B7Jv+cZGg8uH7jGP0PXnA7jsqZa
o2S5oYHPaX4aUvRprMhHedqKBqfnzFu6htRq1UfBOSve7edG5s2DVqUKK5jhEK4nYTbUZXOdMw8T
VpIUKY+AbM9A29PctaDpEQuHf05eeEHOYvv2sbHmONhIfqz53lx5y8QW5nky5FxuU7NTByucwjlG
2AgTfPVvL3u0LUJqjkiUOlgUc9VwDWR1cj00O7FilZTjnBDQIX3jtaGfwAo/7UwYOW3MLyBnc8ZO
CHWypS8lFEXowTcEsCz6x71BgDMA6wfH54NxOO0JWDJd+b3UbWeoz/Ao0m0BXHvpw+Fk56liHsGz
1qK/HCDqFwjgj3aSUzl7Dz3AmNpcwo6qAW3y2n3ucgcenfMivZZrG6eRwf+fkdnH+UOma0b9a/u3
/wG+gmqAC4LKOx4PtFIsl8BloJBUlg4p8fHnFOIWgoeen35EoOlR529e+3NY/++BujjA7XTsLtW+
L8ii6cJB87D9oHWEfZ3rvqhh7lObIvVrrEHXhxml4y9eJ3cRm0aLhuMNnviM6QIoFRhiBpKAP2Tz
0B7qUOTNRDWIqJAvKl74cxth0/JVggeW5SNxpapeY0lUekU0JUxh1RltxD3g3erymXxqF1GKsuZ+
+zVI/mP34nusk6vogNxaVhfGu5OfDXBNTGOEE00rCy2oapIdXC8Go+/aUE4i2eEGPJFi0Rr/WZO+
oQQiThIzqCzaFlb8ueZKfjuVFK3IdMk2loEtitZlxEzMAViCxeOxoChvIMukkLumII/bCuwKKVjF
fGKY83Zg5XlRZ6vEZ+KaUghM6lm4hhm2XlCMUHR9uIcaaO/R+nT5dnrQTiAeG1dJGWKsq25zG4h5
15LmLjmRWZE11m0zu49027dSDDjCMcP01urAToVn0Ry+9yNDYpoOYabMnuPQKrOayOuCkQKNhx0k
IjynCLMS5ecK7SQeDeCkOsJrHC0za0hLxO3jwzIgFYYo2aVEuQc6wzwNrFlJlweuzHoEn5GXb+e+
GXUBM3xRi9aJuW0YEk0LGu+H2eebjzGYkGInbgp/iOn0lNGsJKWwmSnB3rTnJ06XIvBivxgKaJ2m
JL9mPiBuHQq+Uy3karwI1YDXnYusZM61ZdV1etZYaGyRSd7LgM8RvW8M98BiHWA/Zi6c7jSrmIJ+
NuvaUI+aDUi7hkg4Ctsn98gQxjad8g10H1IILIMaAmV57evAnrxWBijZG5MJcofki7Lv7sb9VITX
1j98phGJ9O1S7CWPl/UdFVrSSIjLKU3121ya0L/D6LPxdd9Xg6EM0rdAWMrZ8EkRvIkAiw10sKCV
7KkEzEjqSM5Vj0CxFbAKjPO/fhQooHFmI9ADpyLsH12bynCqQKhR5Yq1WantfKEHM++7pRvRzEt3
/ow/8wRL1FDeapHZY2Tsi6vHDDW9wbZ1UeiGGRUSz0gONvAwDT+8EMjIC6EongLi16fGucs27nKn
XXQ7RrqL/wWRAIJU2Zle7rv7KnXn8DcUTp+zm3pWfA21atX/aKE7x+Q/87yrORs2IziQjmBpV/fe
DkaQhHNXPwQlIV2qkOU19TqJAgJRyhnFjOWgVmCjOge2w8LWQe/oF4Jigp89DUN+l6nH0FbSQ/2j
WcAV6l3fKAkbz/28YRlVbRxLZPRoZpsaNlugA7aKGMtg6uYYx8LmZtlnMLZ+VkSBOcrQIaR4wO9f
xzNS2SU1by0jbgHguDshEPJklTas0p1T6wR7ZfA8fNURiQedrkgN6RgUN/e1X+UANWVVDxtD0WNt
YiyIF1MG8pVLuz7YOVvvGOzhwIPZ8MeQk/TxR/lss7JgLo5v8ljpZlMWXx+RH9aHo5elbt9HICo1
ZXDgEtuoQtF2RPAZYmRHyho6aBzTQj68FJzVN81r4EVIzGVdcshG3NjBsgmKRqslLfC0jGgYVEHm
qh7jLbQJMDeAuH/TnJW9ADxvPuUy89V75awx7CN7DkxaTd7X5oaDYkv+6JoaLp1gf73Svrd5hf1I
DtEaAQDXwBV171hwPXj3CF70hHdlGLxwna9gtmmrwGdglwC984dtegVUH2Ucm5dbWTNbmtrP7sFo
fOcOIiTUeebqCPmtvGpPZlYogk0NBnmuZaSXCJJ3D07c7jYUH+qglbQ9YXyibEu+vqKgcQFE3BP6
8tZn/cnA7slAu/Tw6ABtoTGd0oc4Nwluotqx+ru/RkOFyrDGbNbMSmuAXmHGF7JNpAreF8z3HJdg
yoTQ8Pa30aZJ8ZLKe2CXMNX335DgdfYnbCOvMhRDmYlAcNp2lkn8pHFyrmia2K6ZJZcBk5ZmZffs
gazBOn5/7ufoWxQUYWqd77tX2Ng9JqRKeHFNsdnu025YFjZ5L5dUo7+oXu+qvugz4gfet8sj7ezf
Tm6kuxNqC+4er78FKdBSYEk+HFHww7ITKEJozRMWPfIaNWarFMvRwKWl8fegO/CHyvp4Pa0dfWV4
K5q7zb33dqCVJaDsxvBHcmhfuTKdb/Nw2jG2mHSlQ0K+iUran8RoEeskd9c8hzudhgfAfA+0XRpU
DTwGI+QlIspHPxlt6AXw+7M2ZE9B3YSEZPvj1YbHYzAUtTH3Y3XuuqkSzcLCL3dJmdCDOC7SyCNN
Pyr7u3/yZO4FM9YJ3hCnt7M5yQRZ+I+JTkhHJgMTpb6LBKLnaWggDlHWOezY92maqPUFHyf/SZGS
jnSj9HnG1aWn7+cj4NuVnFEJIHTyTcP/MANyaSml1dZX1tRKx6rxhxkr0U7XQR0Ch8KQl8xIsCXm
Igy6MBGZztkpl9g+m8T/2/lRNWyPsGYcfumeGZRKrvQHlk7cX1HoKJEXGDwyjTQ/qGMlzxCe/uqh
tb/XvfB6Sbv+bbDb9QEmE8dkbv74EvsG43u5FCmQgG14HzZAaqttV4iXmXtyxwTMfDqfMwxkHCto
qXpwhOCrLc75EbrQVdKFPsHKTXW2TCBnGxW2Woq7/aqIHk7mooMKQHSFekpXuXiktzCTnank/wZF
poHzSOCCYiCtZZhpiCf8x8IGQSX9Z56IFykrYzCDxE12kqa3D8HAhrBX+0DRvX10BsmLbmucYMao
kzJez3TdyXmgUbuW8xqsjLPK9bQBJavbj5vXiTGsBFvcaF5L6H/lXi/uwCNktabQ8EN4ggJSCwDe
OzsAVB56NGp1MW58oahvdnsBJZCO9eRRXkhh0Ho9Aw9Ccf9LK4AKoA+Zt2N28rR+3fvr+3d0uMuQ
CH5figdCcEYQAZyHDhxF6N4JbjAxRsSw2l4ddNjqWnl58pl9LC9FkDInAPPKfrn6XJ6xYkuEtEaz
0Xq2/f1LU868wumQbHXaoWgDRmJQsntzOlscSvINaJ5ZXWT2cyG8ZydyQKMNP5SqlGKQoA6ZiSN9
xydQzF4lrHB+DwnDEsss0n0K6fSdCr477cHSV0Wte47D+j0OR4mzbVAeDzUAMzVDzvzyWHN5/9qj
NpT10lUWTvIQnRr1IEASHGh5V9qPlxHq1QQ/9kwhB5/gtu8nATSQchC2hUZa7uFF7bNoYuTLWYwI
lf5SQ7sj/tEJBMNh2RHUa7EB9T6qBoJACsAVSdK/4XBBWIOThXfMQ8BAW2sNYE4z5aRCRWwq8Dh9
iN7+x9pikzC+4PAlq4nltT43OYE1+qdY55Rr5iaXcjLeuD+nc2Fw2W4/t+Ts/3t2HdMug8e8cj2c
szkl8OTdyByEf+9SxsfW/2bhTxN1LaUfhUrrDLgzzfhSGD9RZLDjM3KA13nuKeX+PQVhvUB8m2vL
QrJ8DbiH2sBNRM1hfSnb64hJuvfK1mUxYlChAkniBSC2UqUmecyqAlZk65Yv6BY+axas/7bNkCYV
WCs3/ke89eU3DQyA+1c0A9G3Sn8jAQW2OinSyp8fsNl0M1HyQ3S6otnhgiqgE96x2kVdB25/znUq
rvbLrPq5nsDg5sayWBizg4Y+E+8tqPt8O6BuXuat/HRdb9K9UAop6AT7/874q+/Sq6VcZbIbGHCk
Tj43uYBhcQ3bxH+J9clGqzvtRdqqyMKTpajVS6m5/dR2iFKjP9IXYNf2+QnIb6zNyAPncIyjDd9r
o1sP7gbLpPEsi2q3iqKiJuzs8gBJVTYlQo7Pc4GMvAPSHo1BrB91x4dCeuIthRwSH946mBkOBnlj
fKzFgEVb95drTQtjLxLtbJZEGmmfDphWAvpo7Sao9lCh38t+iNVpTLkXFxolN2ZFY+2azsjCzJ+w
ojELZp6+YC3DMO6gKNd/ZflGrFawynxOEb6CSO039KhEOt5KPvmq/6zoGYt0HixqP3QTXAXmJBdT
HHA7Ybt7NMe8Q5oZFSrsN0WUMj3baLRc7oW4VLgLe2xqJGgPhDHhkk3nAr0pZsKO3/n3vXPnomVv
4qchTq44HM5F7rwLFfmylPR6WNq8Lx//0WnkTne01r9CQuyPV63anTSvXyRUZVbW9HQxLKmGvgKU
ReKoTEKiCnRg+3cl47s8dg99NdFfS1m+goML0BVMqCnaej8Y6qD28N8H45Vpla8tcd9iI73CF6z9
8ZhsK2kHjhR5Dub2tW3YSZtYq++vkOJ590e0qLfYW6fP6DyRf3TDhYkBCaCsU2djphIVToOki0nu
zZDkmiYJNZXsR23lu1utWKcl2hwQlQeCCE90+unhWyVpTq3e31gTRMk4BOoyBc8n3a3p0CMnutQ8
r1iWEa/1KlM48SmJyGMX0+H6x50D3TGz3q4kH1hPIM5U+H9zLovEksmTXQUP2EPPqS7e+jwaC3wL
k5keP6bcvqR8dzO8rfEj6VV4O2RjNUd0NU6wVpJLtUJ3whV13R/ORyoS0Hp++Ae1cq28qUYRosC0
A/3+PT7E3AwLb8ipY9nBXcwsOTFhCItzi3+DtfS5Lx84TAWlpWBbgipzy60hRimj8H1TuDpIEhb1
eRrsd/X+LkkrpfAwsu0h3cYyhbhac4hwgy4rkG36g44ha/a9ZFLZM332BduyGViM8o0+wIhCsSLj
EcbtEceo8UV7/zBC22YH9wEYgw2QuKshhn3YtP+dke1qvbH5rjx8m3FBdioyOZlQh2Ix0wVyiDu7
2lTkVLQbytrOkPOeZ8ZVEzyJ5fSb8hMEMIAXEZDpuJ5KnqJMKRyVI3M748eNtVisKpAT6f4lCcO2
3we7cwoDKytbvMUOSbKAKH0Y2SjFjspNHmhPI0a407FNR0Xs0M333OEQs1unZpzNIQz46rUEf6JS
psCVOvtH+Hb6VRQqKmKoBc/fFtpjZhvs98gPhlWQlcRtngtCBxsvnnSqozxgcxXG0NGKKbANOIkq
DGkgx9z5TFHsXvOz3dJVuiMGfqH/o6RfF1Mn7cWG8EbGDBPtwO7WvznmqNYw4eUqOPyW8KdGjW7P
1FU42wgRJ85PFPx8cekA0EX+n2HTw6Nr5v0r6JBm9ubPb0eDSarPrvmp8n4zg0SVsHbZjBVsWpT9
l8UOsnDvU/QUXQEFAbxmCjCnu44PEHU1XQoZlJi1HBk7HoXkIrqKQ/t49AyF9i9UmqKLCaBjXqIz
qOKfTA6kDq4juiobqudmYF2rTUdD9GXmQCirpuc45kSd7NR3PAQlaspBIrEE+Ca6I5ZC+OgxesMV
R3SnXnr9Xqa+vn31wNRHmXDh7UlmiWDhSbtOvMTqCmCGCrSOc3bI2oYKcMC2OX67VMyC8kjx2/wu
vOUKrQmPMP8PfEKyBNQ26iMIN/xicnm2hptge/sPpVvwg860uIy49vULLa6tRZOuxu0dN11WnUbj
L4j4an5HsmWdBiVu3aKmbtTVLSyhaSHiBVHQyPMx2/Q+wc7W3a5CeyxrCwDUv3wmgmMqOVUYi8hh
UWVvVTUBkrs0B4O5STi7Du46SYLBsOHe+6hYnE8lDYYZfY/RwV0zKa1H01ol6r9dTtMkI/X53wVf
aMWSgvhYEwjK5Us1dhjfYjM/3aa168lti+JOsRNtBGFURqvFwhnm2dCC8y8RPPZybX4UYnuWluw2
TDeuwVxm7/KqlE+PVQtJ411w0jvwr4TjAqo0hyQ1H2J1+QfF2vfTYvO0AbfvdKeQyOCAfGiw/ELU
4drXp5VramoeMcZFEI0coVUzyolldol0P+OuE+72DJUiTpwVZCE7piPyX5hWtWFfVutiopH14FYX
zrIqQx+Pjy1NAlAExI6qxxUjKlTYFbX9GgEVzPq7VAzHyV+sqfXflhoDKePSsBGyxedTL5K1UyqE
bLMy7mfBKU4QWOMTS6acERwRlbLd8PkQhxbKGchBrtkWn8guh9Tp5LQP4Hu5cxAPiVl1xR7S8lNN
FCz+itNRwpzs/9EfW3OnJNoMfnN5asV83HQ4CAGJeb6q4R68ITZNOKjIZr1bNZN9nrOQj2YWGQ6G
urn5EDRLr0GpDajYRsijZlLvxQUKSr8YkCqsj00M9ofSWyM9tSJb3tEVSnivDWYcs1hC/uJ/K0IZ
u4frm5/DCPOesIza9WiaNtRn+1Uf04YvpC2T+eSfGRVgnwCuvKi7IJj5/5AC9gOlfxGBCpn9+aYC
kUf3DW7t8jS78fN8h17W/SFl57+kRocWg/FdRZYy8KZQSymsQsH/Uh4Gy2Bu45Q6n2o0flRbX9Zi
Vi4gOanZ4GnN5hM0XxKhl327a/ChDGhC1Klm4WEwnt4YkaRBiJLn+aW2gQMsWZ3j1DRUAKFQp8hZ
IhpPMetCubWdbdi56sxy1EdaaM0IfinVEwcwuurAME/rIYN7B57cIZgZ3Ih+BU8w8p3OoImtTM6s
S8qTyQzPXYPgIneBNCseMoyJNupKPiUXvnpLVE+YYUby1qs0tiFRl5DT4IBpFJxVMykUuX01RBCa
rU24pk80GGbvwxv8JqqJRFzSJzJMiedmMOys8PWpYInkmJCNtULNqZUmSvd4TJeiyETtdGU0jVPV
R/uz3ZMtpFGyJYjSNsyZBl0SfUtJCe72eyS3VkXBqVxThGkGhgnrUk+6wyLqST/DOJfQLPaUwzwM
NGtLgm2/zSpYRTdoW0FqH82JrNkGhgxhKCsmcS21n6j+annhvYYe3Bx79TtPGcn+7yRccnHHyGln
66ikTDHJ3ii81Tj7BZks+KH1JLU8bXey5hEjPlIxMrKZAiuGkIut8pSZQBzu55QPSqqgYFALQSBR
RswjUtOmD+gNeAqRhUxxQ2dLnDPB1BjNzfqIzPGh0+slrn49gDDKXiREK3MSsDITCO5BNTWrzTAC
ov7ULynYANmv+JGcz2KnuFRYBTpwMGrdHiXQkXVH9SgHS9QDPYij2BicSMEFraPuU3ZbRpMdlWCC
5BTuF0kMqoyD9MXTQMVN6kBEquEy7J7q0wgH1BW+JdjnNL/VJ9lpR5Kjf6KGd83xMGlxn/ocgdiL
hILoOvjypnfU4/8cXR9aaD6B+z7+a5lvFcnn5Xve4pfeRJELf0wQRBQA5ndmBwjLcEtCgGt3YpGX
zw2SNE2sy/s8SNi33CRX4/fw1FPDhGqXmwAUvnhUEtotKY+95KqGTNFkBQIOLHRQrYsFfwnciaP0
I4sjaaE/UeCRbgxcBBof7vpXG5drJlrXGsU2Fq7xuC9BsaD9FvuApx6YFCRlnwR7hzMoVnGS8vzx
r1rIoWWvGmta4VkJ6TqFRkSBXD4FXGUPGnjdc2lZQ8EBHEycGs+wblncJHdUo2/x+j2Rm409ZEPX
H7XWBexRxTpdkN27YiZHC83myqcl/BQF33YsZf0uOtxoVL5dNGa04Rh9xjOvHSdlV8VrLJOB38RP
9FNuf7hBK/XvOJDES085PTLKRUqL2jYaMHhy66liCdzQi6KLXyHEob4JxwmOpLG1ZKdGN5rBlpei
wIqsTYrHDY930gBQM3ucJETPHun/z+Qm6kk0+wNqLfTpfAXsJlPlI8EvYVrW0RAWQmjWc/exaPLZ
fK7DoIAhkmZ2abOUgsmlXw6sHjs8HBSyfl+ZRGNoAG6BHVZlCOmxBM5qymeCyNs27i+Dmlh4bUxk
SSMMcXaapa/Xvxw2goQxc4T3ofTb3ztgZxvoQ6IFtgZdu1ash8VVO7bzDM3o6IE0ZAFr338/QIvs
r/7s+8zFTs2XzJU8AxdwlOHKH8IK+/cvD/ROTPePY8yrnpcjbbA8BzfCZ6djxzLlyiXnzx9dcylM
mXS5szwxrx68aW5bCUT9EuoTc1cz2CjVwev68kSqs04Xch7ZDsE3fsxdpQJzoY3fdB+VuE+mJIWF
c74CVNhhFrjoCKdDvM25JsV+68YUK5xu8IGSRTCUzdfxvkFAGLjysCuZ7Xy20/lDXEKBeZ3DogxZ
7IwW62sRaS02DccBRyUFCyQwMuH6N4UiOCXrVuTzCv1mW5WaTlLk5QOoCBxmlgHHn2ez3bOXHSGB
2MJXEoggOdN/qGa3EZP2Ucc/T4BJbWsXhQ2MSAkKENMgmDacEN3E4l0k14K8ZSEplTaeBjmsqJH6
poWwJRn0RTqLH+ZUXf0C3cFpL6G7l7dT6AzZS4J4YxePcLtXvRCQEojYQcn3Fv3cSvXVM1o/yyN2
KF+FYlQsc8B+JjNyLLTNt/VhSzQbD/eJj8YhQKFxj7/mioVK2q/NPdrPXdTJCHaQviGlxZhFru7+
kN9eJhZo7iHXAAgWx+9IsvWTT7oc8HcEx1woiZObIlpYZwqBanZ2B78vGWXv1joSi1CHPUdzu2O0
FYyz6N6AU9MUiExsA3GaI0w1U2Echh6Vj88XuHzzCWmTzYIEkLZgU6rduQGXNFMv1yVq9ptNjXIJ
pJvhKEGTAHU7FlsBWBuAvKgpbdgQwnCqABd3BWPBMSD4spF0/7Jk/aLYFEOt126ZH2O18UGz6eEf
MB/V6GFUWxpYbg3o19z85H6NNJgGGKwGybiIGCEOpZvzDA10Hz7nEx6ghXqm+HbsPhMxpbxc973s
7naVjPwZBuELTcNcn39pthDqlDRl3Ey046DDEP5NKKFRIXtoOHDA4rOICZsFT80QOIWJAi9KLk+d
+CWuKxwVd396i9+bOGLTqGn6AAmLsk5bmHiS2JtfW9j8DIxIFKslMcGssNA3H8ovaud4K2FkEq69
O1vt9GgQAcQ0D6UG1UnQt2S9y0N9Zo6gESdG/YfnV2S9UwYCpY+AjUjZ43DyG+yfIESzHN5frj11
oJ1qom376aQgKArmSdAYUng1VudjwGQPZnvQVHFfT4uAnrXZHclmN0p0IRaMSOtF5vlMMWFqBVfg
qMfYXKMkF0zStz9YS2N3gY7lXHDLkMSCS8Hh3gnH2hc+OpSoKEDPfdWCSJhMfBAu7KHTachVF2tC
uCUWQcePHcQI/Iyuda1hfRDq8cmc1/MDBX52onN5CoxpRsHTLO+eqI3VlPqimJkOAaEJaPM0PhjK
TnxLTiVC46OREd6avJUsFNzwooBoKtbr1dqEKh5PHRQDXTRA3juRFr2CdcdIu3iJK405yxrQXahl
JZODv4meC71Qu1nwgE5IoLR50ZIzpWqlsX1iOuRE2RUoSRS7JgiSNZ1BMzCh7HeyjnmPWRhH4PC4
LFJvI61uGUuGkvDpra803xxHQeofNIE68cDX7QJE7+xtTe3i1Spnb55uia+WnstOonG35fKIg+s8
r1J1Eq2tJHyBL9wLC+lwLpeioWmC5nEeK2rhSsLabQU1uoCYe1I9QVpllIk3jMMTv4omyEVYmnMB
1tI65T4+2rPrnNJSgoBe+WvNfiNaMY3r534hpNCDhDdnVpvhLm+F+2o2Rl6VLLlSzGzesvSLrB7m
W6+x8GGQfnJICpqHwrbNan5kSYej1STkRAUUzEtUpA/wbHT5/xU066hIz5H8YgdD56n4v/HGaFFl
Igz1LPnKGKzMPQfLwiWaIQTu8YsG2Ddg0QYxwaqeQOOLxhb4VpAaJ5RCA9PNROSEwfgUFOIuyt1x
RnZMyH1UnX06EZQ1pYjgs0AOrRWBpNMEjQ7B0IRXmE7ELacZ61tkZ5cS3KZh0pAJzW+Di1VF7uGS
eWmDp65ni5IEi0eefTjysTF+1WiF0prM6rVsQiYcqzOTq++FlsRqvS9FiVVQAz0N0qSQyNTtv3h+
SwBNPofJdJEzGlQuaYwWOJDHj2SmYH5/94NL3DDUaeBFXcjK5+bBVV8BXlVnZTA9af5LN+uxV0BH
43CQwbzTYmuQsh8ZBjL0BseODa9iG3y7Vbit6mnpggbDsU//Z5FjQ3W/OWV8If/kMbrxXF/Liyqh
XuMfYAkHqHgQ8nYg4T4ZYrMnwvx4V1b+3FpdHHHBoK9q+H4Nz99E9AbnqiUDkAdpkQ5/AGTgUKWe
/lwiYz2kRV1u2SUnnwCm2+c1OoCCZ6Nn6a9yABfnRH26BFaqWZ2SXB//4NVkBsxDmaFjy26+TWpj
czy+winb3jpKKF43Ohy8EdK2GNTrJSPuu8hQKL1uAVDLuTa4cbJHAVr2E0Yqt3MaaJrzqSzVAizR
C1JpJRSdO6DXMCdoxFlPhdMwLeUZ1wa2Q9lB7veAt9nlsVRfe4EAT3hEj3SolDbL9SvctSxa3PX/
g9x8lArIaruEztOmBUgC4GgcWUjZ5FHWt78mlOkiaihAZkhq79awKJIDeRTIrWM9ZVYjoymkcEKD
rJa6QE6hpMMVYvK8z/SAugjpmTZHqX0HkhmC5429qW3859gqZukBj6WwQsk8SWCxrNMpIrtDEOyb
zzsNezKxDX61Po0ofchBR43naS/4HTTnmEdrzG16n6vqS0hP/WZYndpK0uU0MGLLAOG59ETM9qmy
x9ew8S3R524eGOuOFbputR07LTwQ2Tkk6XSKkAffGfH84c7WFQWF7nsuq85xWY2H/9QwEWzyRDEH
Gg8S70zdt0wNBbTs5inFt2ppT3lRDjYBYJptHeEJ0XpuGJWQImD+pZCp1msHxvyRnXGPJlBfDQr7
V9lrBfbOhuHJB3ILIu9ej8/CUq2xE5ZsNQqnRQcURpmDLL8BU4IuuabymHKD7NAh5NY5iXotplzA
VI/CJMv2nh/NMgjoperEUthxa/xtvFojW3h/Ma4FWH570f6kybMXHl6ucqZB9UpiousmphtkGGLu
ggh81p68FRewVaoIBa2tKscVJlzpqURz9nRx/YOSHbMCabCriA8RBR5gOu2SKYA7qZsInd1u+jwo
yCGKLAwXVsLFd6/R4LP2oGDFAX7+FRG0flkq86qPRwGeqa7hpYnyP2q1/G3NxNT7Lk4VhiGfPVZv
HEYVNrzalG38AYdzVivYaiofi7WVo4kC4DLcVMEUmWpnocn8Os/tRpeJY2zOBpbtNRaxRaePWSOR
cP/QsX0YYy7SSBR5XYwcs6TFyiNAzITdwQMdI79MdcCs6fmAvi0c2TtydQ5HaHJb7XcC/W1tEwnj
ksNKy0curvZZ/42EGs5b4gZ7sNAtbRWIPoIyTkJ5R2+1HPoNYb2/c7g2z9A+8YeChXAEhXYPHhGX
FUT+KCGxBTRGgr+8bn/8zco2au659dN+5ND+UPJveE3OMfEjQ2kdQjvZsG/WdWT6+43xl9+NCHC5
Muy7tboU1+EFWriB4hxzHKkayL7meRH2gnbpmYoEEOy6nqd3Bu/BLh6EOEcHcqLsScOe4hxWgBQy
HjbQ2AyIBTKPfq/m/pQILejd4CsFY+zVjYeWdEbW/Ylk2HD1FZZXZ/HgEDXXcRpQ44ZbQOGiOE2W
P227fAlIV6n8nrDNQuoXqVCihR5Hgc6kmAaMz/BlFXbEjEB1LBWoVYpyfKIs0bFJ191/yDJq4HA6
vF/h57rVGPX9EQw1CuGn0Le0AQ7L3ExY5r7gKcz3OXR0HYIdUN4OWgpHlW9laHzh7KwuXTuUHBWv
bDX+s9hmn1bPwIXFshcKrU4k0h4IvuYZpUThelUoWkafgeaB+72YluPRBD6c4V0d7ONpLZlsk51I
cUwdUUS0C8+dGRXr7kYIGXoIPJKHYLEIZypN42YTMqjOtbvru+2tDWJ098G6S+8w7xJ6BJsdsNCp
sJlPrc9I/cfFv5inFMjSPmGPGWf9l5IRU8Wu8tNki8PSvPQ4yxFXyItClzniGqqZHUSA0GS2B8A7
cuUd1wBnVL91DfNR57baUh7F2TomcqQ27Nfta8s8xuowTooFaG2KsPROqJxZ1eI0Cjc0lfo1m58X
Ec64ptjN8xdrRZmnuXMHnu/43EXswNzrTwVErM7jAQxdnvtNNqOg2JXqXiizt7HYtDAUElvvS9hN
R4hzKd8RfaI5+i1VlP+y1p861SWiRwhBZ4yTTHy9QR8RWoSvx7nMBYf8CusJcwuFH6K7SXKs82T/
ONfEpiqSM3jt6RHrKOYWF9C0aYtTvRDyKOK5iqHpfsVDDbMSUoVds1rjifrunMMHxnLkimCbWR1F
rADSMvUboIrwLLNYYQ6AAAQBzzrRuMmExnm8Vp3HHySUL4/H1KrOJiWZXIhvHcS7PjU2JMv8KogR
55ROeOO9CpjNixoeMZfdOg1QLQSwNotY1kG1jSZLTL15R+t0bLQH3U28SIKgJNW6wDL3pAY1sHhf
xs9YUa23K+ALQ3lISFuZ/E5zWXWI3qPvb0lDb7F7p9B2myvSQujZFN+KyrGQ414Zpz7VvygiOVAq
4pTzrBE1mBfaDoqVrKjCnvMBg8QxtUp22+EPZQvwlHBNKCPxpLzFRcJitw5tpBH4uREPxWbZWBZk
3G3aY97B3sGgnIfZSmXVtkTjelfo/1acqMZRS92sYMddyUVZIGza/hFG3P27FZV2ionGua7Qo0+0
crkBwMtG4hvykWpJWHP5pNCrJCr3ysUsop8tEB+ZhI5j6FiraHtqV5w1tM8D/lRJdLJ4rwVBM0Z3
UnV2uu0LMpRJH7URkRRXI4Fu7s17q3wCgxMoTl3Z11UfNUhg6cU1wdWRrzTrpkKa+krdRGAy73UC
pL8bl5LoxVJPtmVRyGLnwRjHLOeOUz33vBMtmYTz59q6jL3uOn7zZMwGzdkE/F7VXEIKauaOSD0O
J8tQzrTxbSK2GYMXo/WFdcNo4qGPBqdDYqmfaQDNtCgSB4/MLootBvdy52SVe2MV/WdFi3xPUzSl
hB58ZK1nW9S2x2x/PPtg+DW2tTAROtrCjJRlY7XXl++hyEFSjXc12j2K4sWNJSoG7dclGaiQM7K0
2jp/VKLlmlTeG21C5hUOB7nlTvSJ8fD2LNFt/spqeglvLv0M2SW/9FAeetxpZfpOQOQ3xugahfzb
rYCvBRO3JivYK9FCeyCGS6ZY4ZRB3WdEHXyjr+55w5CBKTdOUD37QW3kretv7RGyxmXXDfeP0icD
mIYTvwlNtQCfwo68370uWkN3GDLzPLR+G2TkB2Wk9FEJPqiKbOdgOqBa6EW0i68lpgf8s9B4X8ib
QWECjDS/elPIPxyQjjL/tC0C51bMtXz9SASnA2jgmOY98M/4RApJ1qgcBpK37tUTR7ZhYimMNOAC
KOR5FEi6J2xfhor7AOHCwjhoVWxr+7K+gGpCfGmEIaS8Q7oc8S3d2GcXuDpTsAk/6UStN3tlTX0h
BXYWtTnSgR9AsZKug2F2HRQ1N1ic+ewJDBk+cWd30L3SFCf1+DvyRsaeJHQCOJnuChcSn9GOWAzb
mWLOqZ+ICuqNzM02d0bBhb6HvpeIKBqxm8VuLMrAmIxMzeySsIXo1yeL+KlUm1t51+PYDUuOQj5P
VAfpFf7IJel/zFIvp/njf+QGPi5L4RGCjigTDmNoECjgGC9BenQUiZNTcjcQ0vNSP52qqo13kYWM
erLUAs3R7C9xtXyF1srU3MpipAslny3FKdlG3zqQ6tS6++p7/WCnGJ9KGakggIvrEts/O6Kp4gnz
Frbe9FCoCST1C5jYU1+tgJL3x1bhCVRKrlU+4RHgcXmcn4duO9TwZ0yOYbaHt5w3HQRvqv13GWuz
ivVWJVKDmwR0JuNdSPxDI5c8iBZ4TSHv00e9oqYcMDyykJvD4eMME3gYP5TtTNrbAyIY3vXOlWwk
RHCujkC5X4huaUHgdfhUXFfvGhaka7dvDyBfjlrx6d0DOd1KFxf/6dsrML2atQiUsCzaWppuBDv+
AwUXXtOev90FoYtgrNcPtnf388TYvjKc8DNGYdt96Mn3mqF4D/jJcdokd71l8lD+0YXPgWTgG3i3
ANaeIozAmetcsh8S+bvUCZCzD3d5MQFWZh9ChGetkkXQFK49lf34Vx4nZm4UYvRsPrpD9enNcl20
fz23Nwss8AuqwpBeYOEH1rbrLy+qgi49IKsbwn69LyMwCCehGDwSMq0E4/5nr5Am4Q4qu6b9LWIx
7kWclnVmZEE0h7AVs33t3AzU68+0O7du7RfgBqECvZ6MH0t/IZNXq1q2iPzraXgCmeFxCacQbxJ7
aBXpxDd08pz1Gby/2awILQ+lFrWjDfNGs2nj05PSzwYHkfFiRwuZBO5542Ic1gaN45ObaceWt+TO
mFEae4rbvrxS1SMwooTyOhNv4T6GwOwIhAjaT/Rh7EaaorXov7rqyF0ib1tSu00OD+7svnSizgg8
QgeF2H0QtV34LvTNj6mP++I2llcu937gP82dekCCwS5jfmyCsfq1RKRP9RkoKpdeOjgBH57E9Alo
5dcMOn4PzLSHcRSRvUV//e7Kn6Wom5SKWekz6VlbhCn1gHr8vgqHzFvMuBEnNca0eIE+GQhj+xaM
nAktgdjVNeSm8CmSWSOt6+bNzmkszMD13SClDlurE+eMYXCr54dleI5ukjiqiP8R3uNYuJnY4zCm
pXpkPHdNgLiqmxXv6AHICz/fHdZMyh1t/Dj7rBV7TUkljsWpQlt+DbJDhCswK4nhTHh2Fv3+pZPf
zbeJJSugeZ0Ky69s/WYyCJyQDKg/o0mEbTQ3vsngm/b1FZX0y3UvqraRvNPM/4tzZEz6IfCmP0s7
LXpLS6cAF1brsVC8wEqg4MoVPEO2Vi0XcogU7ayguFqE+d7/PH1SFP9+l/AMH5Ps5IrcqN2J0RIr
2RCBkevCeUQGESq80WQ/envcj9k3q3XLkmhQvyx6H30oB9wMHfBDdAAcFTHJgXO1jA1dC1T/fUSN
8kq596/BkFVU5W2b2gl93JUNXvt3Vl+7GW+KxPFI5+ulJgXFwOQ9WQ/qZqYXFEoQPvn0bDwTAGwk
mJ0Uf40LtOcD9b1NRmCLSUJukaSkYv3iuWRMH44X1mDMzYSU8NnD/C0tipKzO7iLyvAddSAYvHoE
gBxF9K/4+ieAWTJwwAyaDFgclUz7aP3bRD1BK5yFHSgoO3sUi4LByRrD30vF98kENuROpSSD5iuu
CWxfpYc6SkMZ8iPwe8V3lYKq2TjLu69M57dXLEKB8KNCnzrts+lyxcJyIQHGFcoqePNgqeo9OAGW
UaKoibhJG5izI5cG5QENxfcAo5Bn+Dfg3wWiFi2slhP/3CjsyWW/wAzX97MomzGJugNOntn5Ze6l
wcqxtzOC1e1QItc8OY2tFAsgKb5trbMKMo4li9cL7kKd8lron1uhqqxXD6fCz0K5TFVmNM+NMAYl
debZNoxYP4FJ7gE9xSSMjVc+uTRurQy2BJ/mlw5Jhw0+FXOqhDpoPpcZ5vpzfmSBeypR3e60LQS7
cYhCxHL11RB1QPn1H6XZcw+yfmtUGgfqfB8bXtFaFVl6AkNpUSX1WbKD4YB8KATxkiRPUt451JWQ
Dv4ULuzp6qF3n5oIJa30O+sKSfsgZAnjwh42mvMF7SwTQtrx3dsFOAdh4HA01VFh1RgjkzEW3PRn
mRBjOsMKwv+LNLupryDXk2NDR07yJl42+p9LzcOTRV2fhmnimoSAnjXaIjOlmcMNVutmQuqzwvyi
+GjF1GksqMfNlxzOIIeH/A8IVEmvZBcYVR4EyJOIFOg86nPxN7WJ/UQgxcFfpMu6evYx+A5bKwcr
6pU3L0C7JH9n+NIyAZ9dRGCrIGJnXOsG9nMK3d9q73Tcm09O4GPu4wASo53FG646lFYZQaIZw4VJ
VQWa8iWnNhjfBFAv6PhaFMbt+4pW3Z93tG4E6wkyYWeVx7BBqfFr3i/krRzGrbGIq1xTuyllZOYr
3jQiWIHG10DLBwpUASjuQLE/poosrIVyu/ajJJwFeIwPYbZ+aWJnEBtbwTcwOKPr0jJx8mmIDG/i
mNZzuWxaE2TBngFco38yOb/nDKw5IOhgeLqPplK0V83Iwvwmbspabns0iPm5ihHmIu4y2sS9m7YN
yUwArBM6r9uWK51W4ScpYhUDuGpqENsybVfzRYDNNkyrDrlkYxJnMgGKha/fLpunpzRP0lm3RAJA
vCWkGJe1arBzXE3LZSq3oj6aSkb66jv+zFEFFgR3WHYfjBdU4rTEVVMMSFyzgzfF4neh3Cupgxsl
t49GjH8WskVTz+3fYINk88B66pkfvm81iA8RwApPZ31uCexVn6EV8v+G0KXR3G3ymiO56zBggIk9
rSmt+R2QZrSy3+9f01kThXX3V1xOuXZjx0NmGEE6FOmmEzVNWi1Sbh3L1IkfwIgONOZJikcbAz5O
LwYdDSDVJEZBw1ScPHLsOFXrklUiV7DtsS+R+TbZXy5MRS8fBXQo441kE3RF/dHYCpeXd6Q2Q0sV
lH+KMncHpIieoDdSL3JS5KYDXx+sJZSp50T9zr6eAHeWy3FHG/ZCdtpecsmCF6WNE5E3e2PJtVNK
9rtUgWo2dj8cMk3hNk6RG9hyT/FVxffeUydINFtN0/oSe15h4y413cHzxYtZis3728e3ECbb+A0o
JukbG4ySHyRSC1EIaa4iLEvHl+cFSkA3p+sWSUjbPbBlmKiN/Lw/NHdjvZpWMeEmZp7FVmB5V2yb
mnDZLyszTos+j9WHzDHOhLIHpOa3r9/b596IVBLUayOiPo1j7GQBybFYItXjW4Sf5BqMMad3hfUs
MFulIjhE4foJ7Rt0fvwbzQfB72GDakfJt2V1yKkBVHULRP7hbU8QI147sbjTc5JANCn0lyJyafS3
3uvJs3nXNaTfHG584NCnGLUzSIP+SGj/1vaFMm6/1AZpoDRcexHXH9TzS7VXAbg0tbWhMXzpzufJ
rJ4v+9BzI53Vy5gYbd6lxb3ZPafe1rCjvF2i8+HWA+x2qyF5bRBFz6mPQ5X/cz3tKHXzxGvyxeCK
t5qaCmDaL2p3f2MopeKP0Ggez6B1A+dc6z3GQrle10uwhYas/fexTg3cRv+wmf0vahvGjq2dpYSP
UxAOJ5FLuLbf4UUzKpvWwfCLIZQ5/fz3qQXi16ytOtBN41S+qySoaqRpYE8+ULDvYpTFt4fG9Z/F
sgE7sFivz6+0Zs6uoU7evFv8xG3nN0DA5/93RPFWQHnSBdYFpLPFn5UU2elGBK1VBbPc3Lb3Szzj
5j9ztPjqjq1NZb7Zaj0Kv0BRYiGB7zBbQkqfJwD5H5PGpP6Vau2WWonjYMWLVw/yDIqZoHfwrprC
gnu0lNYTd5r7FPIGTqcij4wimaPh9oitWl+EgE0Fl5d4Lmn7unBylf3akdZ6ttIc+CyU7oODiW1s
F+UxykP6DrEexSb3ReIiN4gCHqES2CmK+xOl8G+IOKYysQwX6kazt/11gXGchUEcryFeyyAOGSJM
O6mEk4wvy2DW1BnjjWqUVuRWmXF0f5h8lqKQjDmEJQzJxnljT9NeSBtsm56ML8R13sMCFTfiPDsX
FLigjsstwQG+TVLH1vNL8wZG98CXcL08xFIG2CZHL3mXGOgOFfnmACz/TsN/k6YE0PG87jUWekDd
3p1aUfHbor17GijD5s/+LYQW80IshzVWeOUKYhexD1KUNicdb6zELgOFQMrGL0FSDuWzpplSUNI3
L8lBjl1/10mEtmvot/s9+cwd54J/dy0wfcW7pKrgB3ZyN5pCYao/seLq8MQtfWmgxoJdmyyQcYY4
QiXEAGxPRnGdfR1VyuDXmXKNB0kbZZPK6s2/xNmiq66KTXiF8JBGcVM6E5PenUK1oY3CkHNA3vi3
jaykjyVxhR9zTfBvfL6bbTTM/Rf9z7d27cUrh/xmJt9Kk1FIy2OhUS2UaaJ3BjiCiV7rx0qLd5UB
KzIylEhcMuo6rxn+pSzwkVJR6sJYmJ7j5jVmWBJO/7I/BMMr6a0UTB3R1/ghH1ibVNTUHeduj22M
2w41BTccDhALQPtAOz2dzMpJLIArIeRrOLDgbvqk7kJtVUxItCe0lHjJJYGN7kdcfez3DxbcMk+b
zPnPQuFnOkBVRwQvXOR3zQRG7LRN5Tk/QfYAW3wFqeD7TFCk5Oma6bDsNOhdrdSYCMFesHksGqiE
nm1FJ6nPO5OdA9/08190hfdOuwRTSsjK9Fept1ejfbBK49JGvdWaodPHUSbnh/B/YLgbHRyPcblE
KsJE++i5fSlf5Nzig1RrYaBnFvNGoPTrhRBJURK8t0uEEbypG1nLG35h4RKVXZD7G7Dpz20Mmc6C
qvtd3ht27HkSNT1bLmCwOmN8zAVtI/e0oQKH2+twwYwOxFYrl4FZx3UJxIARayu2mspQEDNecKK+
Y67uTYM2ZqYAIEm2X2bwkLi62qLgDG1cXMUDVf5ROUzNEAA1zNbN8vVAuFbgW/PYhgsB0yRmEybc
jlajW1anCb6KBXZzUl4PcVjI+BSC1A8JTzPcCbYosjJOO8qtmFCEl9VyDlrCQ7q9LDxJZgXhxrOz
SMuRHxXeXTKTox4DFkIdVAXcwza2U4EUZctzdHLEkkrAgtPMj6S4M8fic+52jHXu56qndiZnOYl8
+PL/0gvbHc+2DFaL9VcTkUrJR8uY8nE3ja4rFJqSVlAsAhq6FYxo24TGlXkxbUJTYz9QUNuuFN4e
0FUJKR45SAsdxza/VboNswys6XeZSvqS2KEG/VtvFO8Vg3HmpF3xLE6uUVeeIBpWmY73xtZxU9Sq
UqkQq+StDrlm2e3y/KbVrNt4ffS3+ZcZhCgR49o2nM3IzBQTx6UHcCf/N8LksO5602LNsRdsHV1A
i4maVUC9rWwYR7KV2ON5+/4ePpoku9kpD8yTQU6GRuTixuhyPvx9fsnqmFyIUFYry7BW1ZnSZP/g
UpSosUAKjy6HZwcZwYy1DG/8Hvy6+xWqViVagA2WUC8EWZDVf33ZBKm9BYijmQPkNjkbOdDsHGRs
v7vq58L/hETEov1NfpvJkaLT8tl/nfbjLpd15iy+222jX2bHJ5d1ps6G6DhNXmDWrBAHXnIYRQrp
BOrNvEFx2p9iIjSpHE5tGJhh6ZCi++CnpUzHyjwgJW+bJAZM2w2YXm77p47ZItG4Oiir/anIcmFg
BNkfH4jTIAYsCWA9XZiUwWW1BzLncs0zI2Z/W9NnPDjihJZYinu4R+i0H3uve1FixXCG0ZgWtf2h
2eRQhCKJYSWaeLZhqoFQ9paOQr0GdILYiLmPDNL1pQwA3OzfPLp2E564oTnyO0xkHJvghFr8ixLx
4iwpPqIqM5RIQ03q2jhRQC/9sDSnufdwh1k8+kDR2zNlNxKtD/scs2/HksBt3qGu6lfL/lhUgz2L
fsDoVxYofUhS7PxWb7PN0EbGue1ODOZX+Rs76hVAnPeQWPotd48HFi7/K7Zizo33YX92AW7kzyad
7NBDkBrS82kMk3VClCReywHCzjY1+pSu8o4jOnDMYIkFZRCsTwjy410+L/0ZNSHar4eJazyyL37z
xN3rfrQv9sE4T5Vs1sCkZp92ZNIh2Z1Fu5zbK3HNtDT3ycHVrda7qfINq9+s9ZcvlxZDTM4Z7Ha9
VP4ysgJsH8GsToskQfOCmaTS01GeFbrrQgvUkrNzRIPeB83ojoUvrMxVKTHQXq4eiwTT01WY+NRG
6cLpKCKekhKouZ2vWpFCpI7wxpMWnCqAxsieUjNWglb2sCmGC9cfVj2v9kBrEkoTJ38cgMbNQ9vT
8Dtix4NBgNo4vMUBH6TwMl8irH/O0PIDDZtZ4zTPgNRXwWT/9NtilbDvOeAtmk0JZNNvOwBUyhiD
jpSf5mqC3QA9qrf3gyfnuhIABddeuScyPXd4i4EM0shgSYc12kjYs4D5ISKPQ88+v29FYJ24yrzj
AYGCajZI2eC4DLBRh+5ni18SQ6kddMC3+NqkA3bN4UwQBQ7o2sietO/CN4Z1WK0krkS19ko5nGlX
KtPu2iEqz8uz59Tq9ZtXx7kO3SkjQzXcIDcuWoiahNHQOdm+g52RiOp1eobXfgxPGw9ECXpNJmx/
cHOVDrwKsEAKQAWZyKRQRF5WQN281b9p6rDhrV7bsBp50fZ5vg8eEWiK7jkw48YbbwW3+mUa3Gr3
2kRLbXvVl64tTwEyu2Q1N861ilm1MPYY3b2eyimcJ7bgOCbHMl415KjI/MChoOCFzSfPIVD3AqhZ
WJr9Ey9Zi64IRq8Y279lZiv2cycFDXL3zhKjzMu5n5CAlKF9Y/Rs0OblTP9q428vseLYq96gBudy
HkdCGKV+Fx5IT15FcMl8yW66GiexenTsACoTOcZJq8+2DmNPam/Lrk1rD/DykyATJkPztfvYL0n/
GJzS/35JX8j0tHGFrjNsPv6Uj5XxrusQPTrTN78J+8U8tJZwtxXdBxpBchThKeQgMdX008UGxC+P
zu2Pnh4CYEUvQ5lKj6d31HwjcpjDWwiv1lmQ3dT4CEq58lIjCGXXQAWn9SdcsRGvMFY7j4m7igze
7LqaWtdxtYrCyv2lcGxDRh1jhlYMDQU4NhPQeec/gkC+khbb5RA97BIay36m/3G5niHMmcjhs+px
xTM8KNNOvcorkK+QnN1/BZ5YfsC0//xxVy/u/yLPTPgCmyaG5oo7AOqo7ksO0k5onBeyx/+Hk/zc
wbb0zxhV10ujGqqPyAxqdjb0je8N2zP/4nEWeAjZdjfKCqXCq3hChVtvrxCFmrAdxKOofEQDBqsK
lZtHp96NHW2cnzhlSCZeFWvVVqYjoKn3M/LjxXIzgVeriPUw49/zCzWSJuaPZ8aOSTBIWKXwkYys
yPV19AJoWj3EZtk9rDpVg311MqtTVEKpd0nkjaxkaRWmoe7FgbxIyUaGdkkmtBPu460G8u7BwcIj
VZIyJm2EuxA6qOQk9up3HGiy0KCfALdOen9wS8gIIDcdUXEzcDAJAKuhoxxw6r4KYs+8az8CRsXF
d5bDgz6q/m867vIE2ey0Yyp2svRZLOIUqQ3y9C+2AU0logQA8CaiXleGqalXVvt11VfALgCA3AeD
HeExnkDjPUAhX7hRqvS304H0cXbY28HfwkNTG1Vn7kKJqCDaJ2YTqBnzHY0LPYcyS0+GtsqrykIL
kmDeTGqHAn00myt+PvJ7CgVYUj5ta8w3dYnh2l9wx7GTF+x3Ed8X15TV9YnNarVxZnYJfJeaE/9+
igSXw0Tui4TrXzotAp0iPk02VXjPSpwfSvqY+y7ACIBbyjVZizDqO7ie1wid4v26ehyBJa1c5yLt
h3dJJFGkAvrgA0dRCsb5y4fNDQnpERyIttDsL1rQaQzgRXTg6HBDXBXO5gGRV+D/YwwdAAtbF7y5
cO+zQF9wHdK1ZWocz16mWT8Up9MBF2QFgCly0vhlD8nfl7ZlbtG2CA6ZRN5Vl+vjjevjmSWUkkeC
TW7pU/DopWWV1KgM7FgHLP+0ce/Fp6Jd7tPOPA4+b//xwz58jCxVaE0UEVR7LOX+wxLaK/v4DpLm
+jladsUm8L2TNxHYpm8NK8o6q76WxtHWSCTWDiVDgu3yXhvZAiALiHInkbWcgVE4BIKYKdx4UQ39
CQBf5o0zy7Kx2mDRp0A+h0PNBtZadqx/dWEZfGoT+fzU0YGYJHBZvUWsb2LDXw745TaM/EPjg8aW
9A54qjzGygWo7yXNsTXjcpV3z3W0IAgPlJF9ikyaDXccOcuCOF3Rr9ul2AFdxsOPn1OUvDFbGLSJ
l5Bkx1AG3ixfEpsP1CfYoMNWi2QUDDVW0KyWvcH3vmMQMSHOuSIauj+9ELsoYtOA1hIA4wdJbYUX
0BBDhB/3paoYX69XVFkfhVkomq8EmKclsppYHaPHEwMTw6hQerNya7HDSzID/h8CNoM9UG8dxDPf
3FyFLF+O47leWdxwExB80ONpCsLPhDpepwnN1BAmtOcU45xmjBqLk9iQaaCvxOOS6w9deSAr4czu
sNWedEWaZ3+0bGcL04pHa5qS9zwUQSyhau3qrPTADcYoXyEmmo2WU5sD6S4qP70Zvt3NmzQ2lA14
OvYXJZPnnkEXGtIUbLSP78AYYdjHkHlj5Ea/OtiS/KcmZtFkybF509VZ63V3XLxxGLwlaBUbnVYv
G4rFzKrpRL8Wiaa4a/vXUCDKURLEgEX1EOix7M/218Sq3xIDwSaw5UjAXP3rfjvKneKVVxyLzU+F
MdjesRNnFG6xlJDh1Im2Rb/4WKnGkvDoMd+Cw18rNPYwUJZWxOoXU7nPbgR9oSEEDuP7ROULjrGb
xL8In9iYxYWi8Wfgwf2yTV5zRK2O7Jk0XKh1CQUAZHyofYLppYp3kqyBNOPq73zK+J6T++AmFFHY
gG0qtybR7pos9VWUj9qHPdh+42+dPM6o/oANZOBTHNqzhBlBbvN2DoLF3DHbrPwkgp7oKcawSPDz
QynUARVeFu2D3fTlwhdE/5kI1PYL5bBHoZEdUjv2jGY3XhQwwZTo+JbTSISpW7q+2Ll8Llf3s+c4
wTip6ahVUUj8InvVti/7hxGp1LfipC7hhQNvLN/Mbx5nE7dsD/bWeL0wLV3adzvFGUNqQIGcoVCn
jnNChXYjEAsVziBE65LxU1t4x1U5gIUYkWMKLaoitG+B7lFuOKT9Lh5yoYRI9u1ymjlMFMFkPfmt
TZY12zf05ai8DVPiCDylaVH30qNTb/Wa8LtemdTz2MfEYX4uZy2F9qUbXlonqKQRKXe16abnBomq
tH5jyGe3cU9SVK0bBwNVOacoTrYAcRIBTiyUj5reOPSP0TAKiwzP3rEQrywjjzi1v56tRhjNL7in
oIZfIGen5uxs/maOY5nSDj4eujFpA36UKzd4ZH2QTc/aeqgedCl/OXaS8nPWz+TZgBh9VbaYMOHu
iul4T/MsEsGYflnSqAlIJHkGeS+ncwUjX1CeFXwMHNcWJl+hwKwfY2gUIIxgJTjCfJR3uCs3hcLU
WtMqk8X3Lp5c9NzX0/x5WyH0YVF+IrjRpXQrfEKthOZt7ctxM+43stPhg/Ep8jb33jUUpc3cml8O
LxRumFji54ZjT9RuXd2WedtxQFAQZaGUOTTQMQuI82HB437s/HDQRH3jq4enNTzdnFQgE/BoKc0f
hYyH9HOKThvlndKedFHxNawFMY6eYz3ZIEWIt+rGC6qEmU1MJbnDKwev0K+F9yTiWCNr237puu81
m/PUQtwTjUWlAFzkP5aOWlQNfdMKJbqVbbMRSJac6geI/lbS5czAXHAIrR3thZ/xJw7ehab0Fxet
ovs2gsOxZqkEgHrWS6lbIn3HP10myvmQT3r5rR1m+lChvnbiCgrM+I7qSWiU9MGxAJkIP5auMTxT
C375l8V16nGJtcenyE7HnJrtK4KgOK2UpGbVE+cEDZ9Aw6Lv1BkQUFRAecGqK2psb1fo0Yew61JE
RXior3aD+5qxr+i/EYeemBO1K90A2EYPjpVobmx0OtFejMbFytTEQ3cClJOJAuzo603pTc+WbBYu
3+O0arcdSK7Ltm8Aq1nerG4gQ7VT1TAD5lz/k1bYbVSFukAAQ16RmzpDFIUkshUsRZ6e7KxGS/hH
ug/4uG7DIdpaBEWQSo3Xk+YDtXR/PASI7RSQy4lmmHbowZqggLpido3gFWGYj3GsePBTWRbUtFN2
qx/Fd/+0VSa7QOi0UXLw/SLlhJfPjXh9h0eWBkUFk9tYBk7XLPcCj52U2mLN8UNz1BYHQ7zQEf0O
VM2b/nRtTzQyyNLw1NqRuX26w6Nho8eNp1ghLmuTRHrqc1l8jCseYS0aIpOAvma8i9Qo9tJHqtsu
1tT2C646+UehP7UouhNcL2g0gnZpxxFK+/zBqd3gKnfJLMsek3fgJiiS/Nmznw5sG56+27cksqbP
pykqNn3REB++iPkR1Z/3aJeMI5W24MNkXu9KZA9s6HmoO8BuuchhQEYsJ5reJ8HV5AvfWq/XzWPI
6B52BgTsCMhbi9p6sS/gzyhj+m2utWT3L8W653vGaIScZiCK7GOfaX+0bj3+1KIWVvJiyFi1H1Kt
RCUAHJPTy07r9sKSA8+hx4JmkADPyJcUErUzhgoUHD+25GtzomH1aB+IDp849jP7CdahsG+CmW6+
bMFbqceM1Bu+koAPXuGNjbk7HDcaTuG/f9Lt1JXkZDjrFJZ5csW4Oh7Jjbk9GRVQCJp7uS92DHva
ndgWYwvYUsRYb731L8e4b5jPbSn6im87HJffCLR6mrSpSPguRvlHhTCk0ceXGdtQjjtrpUhIJm/V
GyLAZyTWKCDbLkET1S23gedf0ijr5MTx8IueXMiDMrpqfOgQU5ucWn+yaJXXopsma/kVgUdv2T5s
qrWELQKzbeHzVmCHU949H7KFjVNDoCxslHtIgSrERYiTajzqiLtDdqStOrFVPHbNonbD/LozJxOg
CnVh7XWIEY+8eseoL0GgTeY0s6oOKYzCStFRyKBPbcJ/NyyIoCqylGhDal4DAL8WN8J5NnWBvU8f
1gSFyR0glR1E8NGs+PMKVrFGBrHSdKQiTB+Ft/vViHwTITctRat5vTaTnv2DqWC5uRTBTxtR/lQj
XLlbQj0rpHyk7O5fYmndsJAu/gxDQ2naPUqFj1kN908Ay9T11wRJ3H2iYXIDk6Vsw3eG6b6N0zgc
6/O9334hMowcx0bbrCgVdqDmSNR54f9zRL0SN8RE+FCSnqh8o7nzdywyDdJG16CIe4w8XLa12fxk
+yZCXwp3dqWuktHtRxopx2hla8EShx6ajVR71eprwoICgbKjWT9FTl0koBfuRHygaKlMg+4XpwXK
8OzCQKWePtl6cxdSaANiaUw0KkDJGEhF9I/QnY9eEayyBp9T09ukIEGGKkF2/AXQDhR9bYeXLMlH
FAx6UMGQ2x/98HHyasL+5w8TnMnOp2UbH9Ulf2emFKiKWA9gYicynZSkXxJrqYJIvdUqWyMZmqvZ
/TsQG+WP5XQX0OgxzrT4Tn1DwTGY135w7RhK5BBg34fdx/zzsUg54Bd5mI1t4FsySJ2wUErbnOhs
hDt1D3xbrdaW+vUPM0i8Eb+oehksjZA0rr51NmjrCOYVvV+avzrEOatqNHhGJ6+2JCLOPKqWxbti
+5X0FcLvTwzx6z3mLzIvk/ym7WL0G2vdVnKxmbjUkoVPF3VBOmPRkktdcgvGSBGUwvqdGLzfz740
qGsLJM/1OZRL/hew8XWR2xyO5s/JKcJF334WQ1uPFT01m0hdhQlT/45aURmqpjmS2/iQUci96Dgt
98XmweKPIkaYNj5Ayh6FAJ4D8YoFcy9VIViz/8WpkB0HM4oH4WrpFfO7immPtAmWhnrHhdtm+k3i
0o/iMw1ncErRLPb+RYRRgCjWYXrgQ1uaGfApYLsKHaQ60yKAV11SgCdtx3bk3hcHEPfwk9nCLMym
SiPdH1sNix75oQxh87UdXSMxZOOKdMdWh+vpMtA2+CO68AHq31OxlKvJv/W+zAa7w7mdKI/QKSD8
KrEFDMZT1YF0PWcV8B3KLl0B+df39xEtiuEXGKGK3qO40dnAXk1vjRX99BNijVfP8WlcJnUZfa30
mRgwPqtoN8bzLDbZVmvdIKnzERtebFj3hCWpyg3iTjb82scYOQ5OcTv3ma0N7RCprmbQJTDYCLUB
2joFs7zY99gKi3LSur/emxPdNPq+dBnrlpKHAMTTwsh0jUELtfyIladf0FhCKsOtkg6fsWwd/SJk
Lc55asZE+LZ/OkAtb5G3xZ0hb1hoVf/MBdl7TP8maN0HRwnNmwGVKIMyuuNzifgylB3FXHropOI7
aukXkdpoNPijZb2xOhD27g5kRhdDO/fiPLO9Dfv0Zm0jvsQNIvGvQr1WSoVaJtdhhtNsuQumL+Eg
wKdwjyxUSx52ek16LHLJoJh7PcdbbsOJm3mk8Dwr4/71ttTOQ1zVlg+ygUI0Svf8cTG8CWLXR5tX
62E+ZA2DMvINoJt1vPalpBCSFNrOKMUBrqsr6zsa/T3uoM79Ru1yCBEJGvEB9VGR5iWJRxJteMfe
OY5hpPtla8YWOUEV/a0M8fuFctv34T0ZMuyJdaNGREzz8QQYPMWrT8AUHyDy0fWplH/g3udy0Qs0
OlhLPaYfvQQT/FdiGqW3Y9hBBH3YJRObyOaFUvU9W/Bdhy5U0vTFY799VPpH6xZgZAJP2PPFV9hu
Ovjjnl1mE4DeLF4gssIkSnG/474OY/bb6N971jNW5+CWE6xDe4XxbqidIqrY3IgXGKm5lsf4SRUM
ckcx6vYH5zT75x5QGgb0itlqJ92QYfzB1vfoXUn8pw72Z3Esr8nq124AybK+ILHXO6+u/7AA1CNo
UbhaLaaCkCppoE7mzwnd9PNJeOXjsKBLuETkIKANVBqub08ywfiGsN152Hme5Z8LuqIXEMNwhA5h
xW1JNe8cVYHeEsI6sxv2w/qrnhL1yxfS3GibLuESJXCW5C2XCeJpc8f8tFEbaJYDKbeSoyludblI
tAd5cmbB0bLOEXuldKviD1BbpNjYbiN/YBNLRq0oItPshUDHebx4nCGSsPFCMSkm/XTlRHCEAqYS
0P0BXKccz7m7HXLBm2T62NzaZ8CC9/AtdXk0VjjvBvksHUzuXvx0EMPPmFfl6gm/Hq/7zGbPaSX9
NcVdVpVHTDzgfOrbQ1dei6VfyJ+Uyg/kScvpfl1jSQaBmmZ6+Y6Bz8X8FbnOdFmP8X2eoxaYTHxU
9TmkOl2m0bVQ0as0uYDYDIJ6eCTJB4Yc3b+aQZIbFHCjs3SPFTS17oruZ2Nc/SYtiy7cPNbkFSp7
ObuEgPnI4rh0qTsPyn0vBmWtal4SKm8ZKEFFhW6ZeU1UPDr9mMmDCem1hk4bOh9wareHMHPpXywc
vPWoum8To8g0N2bmODypGMY4TsKMj5B6Sdxx+c2FA6qmRX61fny/WcQkf1ocW07atqU8PZ8gIuD8
rkYxOTdfa4iY9PYS4iZvEy0B14SMdW9XzxpFyJpQprSz0ULTs1zeLvkk9en4Tze07q8+dD8R2gKN
1EkwXskBdd7ag0YqBtTx6fpFWDJTUEXFB9Twy3tPwKyeO1qJ5Iuw7Hp3h7MyzdPOKBi54CclYWft
k+6FbnMR+J4tpX8UGTKvP83BmV8QaSriG2+htvyvy2yKx1fEiMEZ6SkYomvExgYlK4j5gG3qOyNR
wlJH90kdrEBmTTjH/6psLIGAOi9FzIRKKLmVfTo2VYsqXHLrj2eDOP9j/C9p5kVLPBLOksGpT7NF
RInXFrqyxY7rBbh0rpwkoMVLaydFFIKA8ELIcLjlUjMxd9h3DZXSYZF5pukHmrcUiOOmGxNI3eAb
j04F8/aPOWs2cJPA+tbQpUm1CJTgGkn3rS7J9AVyKhQEYlwIjOu0qgWVldgV3ckBTbMNw9+8/ArA
J8eJP2NKgnRR1EWRGQ/pGJrvJ8/ilvjWynVU4hcMTfiDlaSiDQB3ndgpsW8UoS7E/U7BovgNj56I
C/wbbqZzH+s9SXABvGsxWUGPileTc3TW9YuLPcf2z8FKSE7nt1yiDSN81Msr13bTQCgXEKgUViPG
igfUFe0K9pPMvm1AKDeoeV5a+FLH9DBUv5gLXdxrSUt1TZ7+A7rsFErC/AwV5vThA862pq2v8pTs
YjgY+FDR8D58YiK9YbCfFk8KJGC0vJua/8ZzZNblkne49DQof9upsPp9tSjjDTMOpwZaJH3D+7u5
VbUA2x+ba2Sci+2tfPtw4Ic3b0dwBeV3k7ykGsLp6WARWLVdSi1zlwMp5CHUJbeo8sTK1GOv3ou2
azXZnt9oOa1eajYkjwSBIKQIn5f+QbiOpp4GHSXHq/JcgMcfcEBIRmRN1Zg/+sFbU9NY1LA6zcJv
1rcIuw8ZnfKkd+Xair9OHxafBDs59icDXZ6M7exYdl+9sEsXw2WXIhNY2k0+uZaWixc8qXyJCE4/
GhZD8DmdTYHMG/VnSdeDKbKWKHg8UXv3Rsz+VbR1UE+ZMNDIgTyDfduRCbNDiTkEgxX10iYT58sM
KDOLa1HquYigUYTJKcUkxY03uwnaPmfkwp9SIWB2s2pfvXiduDMBLAw6VdqFW/q9NS5HYHuqZO0V
Z+1joPxUq/efu6GpHw83TfVl1hKuKNZ/esvX3yoXQGSKIshcoCbBT2D73Ymp+TSVrV1iRqfCjI7B
V0VLC2bglC9mp3OHAL2snOewjAFb3vd+pZcdRifiZHnymXmU8vNsuOLMXt+IUdLLkU4Iq/jloM+A
cTv1splc6BXUvR6fZ/G1+AlMiMO0PnQR++BTA9CGRYJUIKoKpLrMwW3rfw5mSXTmtqTUz9lwYqih
ZDs54v1z6Tlm3vxy4MYqPGy0eGH277et3XgnwqHRuS8FL9DDiDFT4mZZCSJ5Kt2/tH6trgQf3pSF
OHem9GuHeL67KnAfvni/CQdpryJhgBg2pADQ2yhMx0evi+c46KT4rMQ3Biw2P72kmHLh4qq/RIIR
aGrjutcWul3xG6TPkQHdG/o2BlZ12TOM+bVAm3h9GSNKo3LIRMKkGrcStfeY9BtZITv8gOJ5sctm
9+7FN6KhOoQxIrGllXJWW1eqx79xFQv1/efl4YgHLZhT8qOjioL+Zhh8IAIQiML2ceHMahfEC3Og
wjKIhbkQOmMkppVLoiCLZeYkUW8ffFYLOiw8yVXREvbJZK6oNqjUAHBBrJwggUhvTKbnGoRqDjJJ
GJW46yjkrsNg3y62seh7Wa8+9lRqbI0gp+S8zUkEiOmw6OGkoT69TasNYUcGMtnUHtNw5nPJQrZB
CuEOGin2fjt2vYwKuP5jYjIWpKL4JsYyRGCUQLOp/tyO03kssdnVY1MuIhS3oHRuqMiylWZJM0ig
tJ5kLWXevGBye8j9yYT+evC9LsZoqFL2Kg9va57G88qNHRcaMvJVCoUk6pWeR7L3GEEG7lfSN6W7
yqoNRCe01EUg4CeoujdY3zUDyQsRzG3fhss5iMnQTZNd0Pa3AdAxThN7xQX65SAOCr4Lkw1c6tfs
pIz5xNvI84AMLmlbHSDFJDNu+jsfvtk7NLfwytbCPlHDsAsYdU+f9pDHu+Lrm2RQ36LUXniCJbKh
8hBBbySr8g9XHY8CsPO3zHjhhqRfbChqorvc/G1w7AFnRMZppLG6IcAHAHKhhdHVlvQMWOr8kZdu
OFqf2grwjBmvwCO7DjXBUnUSbBtiNgEkW9nVSRNMZ+qVUDVrwUyM7IkteVPDQfMMfdfo1TuOyePm
Fig3fxsdTLiHEWZU3iNqZuvwehtNeRbFQMzjUwQte8shwx9e3m7/AaS6DIVk3BsIGvYvCqkb+tFT
cdUwdmo/FSHheCn69gHJ/WmGFisM2Icv6zyz9yAvYRKUNDCReIAbmRMBhET/eu+gQ8wg8IxJGojW
CurwO0coCvWhOTFcUk9dAE4/dqbmNi92IBFXrmqDVG1aB7z2/upoT3ZHHDWPyKEP7+xyNjKUfGf/
j149JqwWnLouA75/N0uDtwj6SKq3w1SgNiWcrnZziIob/D6n7tV9zGxPOD5ampz4P03uI1CNqdq4
wOO6fuKAz9J1hXV1Dg+uVfjuGNHcjEgCE7usXAdUOKGLiUuB1irHGintWp558M9yja6TaUlo87Fv
ZoUHkafUB1ppH9cMutch6FZoQM7aCi48dWJMHYq4EyZCDV33/iU8ZjO3PpYbuwUntHhAuqXMgXAL
ZqRzc9Mmow0ZEg7QquPRTZM34DlJH8HXUCgfcVtdlVQt7q6aHNHGxl5cE8s/l++YX698Lg+cgbU5
NIYB+YihHVXHzpUt0FY7WJIRmAQtLLTqYU1T+wRIEpDi7gpfQ+7g/wHeOEsDdXbjHQRhBFjmKK4u
UTLdbT2NaVzsLdkDQ37oCeJ+/tjvhkW3G9ZFs6oFhXTmTSDu0NE9D0jQt77pUwrOojLKZrRyGwNb
RuK4t9hLLoHAyYD7nT5AD5kcskL0pnn9T1NS/ERhUr0ha09g1Kri/gqnSDbkcZUynE6H1SFPe/OW
Rq3T57bFK/stQuMpS31L588Q5QfhSrWao4DWxM1+jqSKGRU9noqntAvNin2jVNQltem2ViGUq1x5
gBqawHhs3ldeUCcJoWpT7Yg7t+tL++ss0JWZucXXNdDMkkGGJd6OXYLGN7CROXLqFn6ubsFgwxSn
OI77F9vKBVSuQBfoGqq2M/o26dzj7o1qyP4lHr2TPIDph+wRLbgZVSo+rRcpUqFfwef/ewyyvzHX
lYzD94GdpKn1gZ6Ej9tlsIHFa54Cb8BEyr3Zsy7aeUA1cvIYPAR8BPxuTW/VtX2s7+SS20JjuvOY
kd+yj2jb7XLJzLUdC3RgHkPdhZMtjj2T53KihLz9UC0COWcaSKMu3vsQbU4FrNzPSElouEZKI/QA
q6sAikHD2ZlRmJIU/zxk+ubP/dINM/kwkjBD+NDXtR0sjezKCz2AD8VZR1AWBX9g+VxkrIybU4PR
bIDeoCgxJ16ERx+pMl4LP8ShFAryc8gmxnfPWS5jaXkO5W4GO3otOhNyuVyBU4jJlJrcPZWGKe9m
YWvCDMOf8ipt+WPbMV7x/qyx4UJLmbOnkvHD2Xruc9ZJPBLln400z6/IXhXUvddRqSz4EXQZvXPo
rhaavYCCCN+wOa2sgfH5yELMZWepBONBHGMufIo7LQdC+RtR0DT/urbq8XjdnPERRbvhDpTpKEkk
1UX42tyAohl6FCEx9mf6JidcaGGfp3QEnEse1rDbt1c9OfbgkDJwii9ksAY3m/VDaGZdMx1HTRrL
LyNVtvq5q/ts6grizNgIV8jDNmAU8vI5/hxkWNu3+M1hEfnb2Zdgw4eMCeaD0h0voR7f2/hexB9g
dgW1dC7X3bwf8m4ghslFvy2ZgsLQQYcjX/pOwYhIYqzdkTWHFNUh5WWeRfmjLEo1xhKyaF0fDxX0
6MrYophvQQ3sjl8NOsJ4QLt6+0f4dTjZ3ZLFOj3tGhR4gXb8DvDHFvrdrhMyo7glefhpXKpELX7b
SjI/RTH8ohf3ZQlhGr8cNCx4SLJk3d76tBGWtHZfVwu1KLa8j3DFsnSXxPV5dNqYso1Jm6VmXhQj
OFzkbEMqfVKMd621vEfflAcD70X98kt7ll6G6XWLB/p/Zix8OQuCCe2J2GD+BgZhPgtsRSn+xU71
/oQI5sQ7vNWUq3fNpnYuY+8lOJoz7wIbtrCJEjKV8QXUQwXcyWQgOWrjQ6Li6rzRjS/mt8c4buKj
f3ho8JXzJPcMw/xLC7rnxgYmxHFk5YKekw45CQBCP82e4h7R25kbOxTMIq9gITD7DeTJ10SAV1TT
Hm7kayMBuSCwDtkP+4fVq5jL9tOV4yo8Nqlw6PEmg+6UwgYlL36iwn7AThPCKMp7s16OB6R3oJ9c
tOOOJ2fFq/HyfUfdnwkuX3qayAUDM9CMljoFKsYXNtHbKoGMA3rjiES1yF9Z9qoS+03MDYBiQxQu
qlilsP8x3F6RjOBip62ZvybdOR0GCtg3VcMhsZMvy1NGnDqjqcmu/CJxVRuXarx+abv6jL2QqInO
t9G7uHdnP/W7eWAXZca24jv6eRvt9dFWFBT1l9C3z/Hx5X1ORrC6Y0eOs09GoAYvC/ZlTfwe2IKZ
N0ilCtKCZT8cb1KWAiJ7rlJBI8Z193a4RSlvQEOS/RNid33u7snDvakiVa1PGYVTiHLIUXjBC9tN
MGVGr53B4okVmfzKgdbYIgjNPUYkHKrrEUC3TyQj5HZPBLz2JC7ECE+hIgEMYd29xlghKIR1notP
SGIcJ/E46ym5n84k4JUbJpzEvl4mhhJUOMXPjsZKGesmdSCKxOrdv36/uZfur8krboI3H0CJyZ8B
KQDzh/8jkqldVWfFiwaZi1KHTDwdYUOL8LgDI3+/vYWz1G8VC7djNK8vvmItgCM2dK8DJDKUUgkM
h365lMpXMN1/L36Jq1vgf2ecDbimRfYxAdvDJJYGtvQwq0yTGNLHMcTWUDYeoO7sF8zYxuUHMsne
KqATPyTRjM7DjmwLFfbHK3Jtq6cxVOqHyRf4C4n6DuMeH3dcwqHc/oGTootBgmDT826FKTuGcqI4
A8ANtwI4Y/UyCyDkHPFwcKqw5QU+8udRbejC5MfnbjOZtC0hBcc0HyZXi9CGLUbOMmRP+ikPhRiB
wg15l7vul6EPSVtNeTNT2WYHXW19NvCi6rXiOTSUc0A5xD9AdafxU5TQ6uH4OIpDJNzpBW7Xmw+d
Ee64Dpzsvgu2rBwjfaM1P572tBSQq7Xj0o2s2CeNOAGkmAGbcxlRnvbp438twc9gSRSI27GWIrMT
MISWJUShVXq39haGQr5DJkU+TOpUdcCeHg56zLUeCbj+1XghsiDp6d4h2yJQmtjIQpvH3gOdVkl7
zy8SHEHtB10gro+4R6uh+WOCvfNFZna0eyGmXBhHTah1G9F8p/q0qlnTFWGcdRDAxtWQXgG+rV4o
V8xQ/Z86GXTnnzH6dXj5DeKJdap/MUBkdqe/hGxPkTG00S6RDwaLgikQXndKndXoq6cmp1TIJ1V+
2AJCY/2mEwZe8NvR3X4qzvZ5vRS7zMWEy4BHxc8m6S6hL5wsBdWoYsUQEkCHjO3lGfAMbIMVzGqn
sAXuwD1KQmEKb2yBqE8aLjiSPKUnczk+TjcBFV/nbV86ZNRdOTpe9mb6Mx4R2hVkyajqaGgqvjJq
FYI2Q1NPW+KrTSW8mEHyenej81rDBFs7qGVg8CL5f0usoOd8ehcscEDKEToKgJ992UR+CHxM9U9V
dGv1t1Jww7srLmCOfJN8EYlZvQ6/I2crFS8dg0Gty9RsKK2RhGmy/jErhHyPoCzSysmchrMQmvJV
1S7puUQG2Gaf2nH1ns92jWNcgwc71BaFpfqVBwDIjE1oyC8dBcy8wt029ixN+xJpU7lb7+tdJUsn
A/MZcjpW2gY5Ze0WLnDlE+xpladyVW+Cys2QlS0+BmTJ8hM+0yAYsPEaJjVMvjKOIogXd/1XsC+2
Y7BrpHnNV6puGWmMu5Z4HKu0vIhKk3lGzaTeTS7ujW/9aZcXgLPCIs2dQdWJQBS6eXQ61c25iP10
23jjusdf/ndjPqc/zCjpxnrefoUszIs23j0p2lrUgawSrJuTah2JGJvddJH8IEoBnIui6k93ejbV
WzeFZjFeq42TrN+1HLBVQNIShPp6vyf+njISgfWUl6og34f28yggr0PWBvoKkUlr2qm0ewj5ohKn
+gahrvB9Fu+H0anBF4ZeEKbH1l+/G8Dm7FVhUeoGvpu2G6iNVcBTD7v+Yf3bV1CzP07j5U0sNqvj
QSc8LZrCBFCTmaFhvKBhjo0iuNs//nSV4r4ARYoNNYW+o/3yngSgjZqdMUBo6SALR4Nvn2aTb4Bx
0ygMmdE6GO5c2MR2KJ7NaI0GCjTvzd6+SR1voHN5mjfOWbF6ZSUgGHQiISBv5xwYCNdGfYA1FSUc
m1bq7sxgENdvXUVTScep5eNmu6cI7cY/M7NUpjqFWvtgJMzli5WSTKn81Fe4tuv1YamB8pljIsdE
sxdFhrFftMO1FB/trbBbg9tZkNGJEyjeuhQvIdioU7RDZhU5WnOgfIbC071YPT/FE8g3fUVKNO9m
83Wg/xLM1mrbpBV7h3W60w3MASKl/iHmO/ItjVy0fAGVmrTSS5b285URgfBVjXxa/JRYIz1uEe82
T3j2S1py8l6svtRbTLapLkhFsYpsT6wwpB1fEh0yrMj1I0+BCW2cG32i75kI9xTYtIHkSieRArwi
8aXtdiWGCe2frW21kWAgkN7ARCPEK6MgbPKW46s7JwKU0WuWVmbaDpnMjdRencX2Oqj+Jma3e6pf
euyS5C8H4rhVfMC1TOCIOsvdBY5CSVPWb+zitxo9e3QuJ5ACIb/gKGp5+FPdzFV8vS/ho2i+5L1+
6BnrB/FzaIKKeS4R2Bp4LJbtRbJKQrOS91qDYJtxD6OWF+GZ0Nz/A16w/cS6arD+6POJ//Otkv1W
JdsIZAVF3YJflz3gYfhPiI0zdRvXApTwg2sVgzUlYqPRB4965jEeIETgWVG8JhBeFGVN/Bjq8HC+
ngJzgHCZOBXFscfpwwo8kPBEeJYdHZ3SLJvRqVnRXpyEWXRIJkTFLIM5fNPfT02z8GAZLN/+DBkb
TctD4nsftsl54df6/VxaKRdV445aW2agDtRvZI4E+r3oiVjHwS5y8CUpmquDe24YvOnoJCEdrPxe
BKrQOW5z/kyHfjUooeW+ZsLRstq5je5UPO4iSmXEi08LHoRkhGublg6L18uwbfnnFn9QjTEiN/eW
SRsRjWCjm0mFU1eFh9BXHiILGaxpUJItk31yxZNGgXhsbU6akvMyPQjGlI72alqbzX88z1drOOrj
jURQhP2UNAfSDeZ5TE7/zAY2M+bdmMjy1wbTqg6kBRQKY1S2kPs2n/nCnnLa6bAs+83jS8g+nSDD
ubBgQBA/jazK8RdQ6FeQJZOHTKrB8S3nySNduTT85IZAwLx7LanJZufoT4dslsxIhiPxvkZT1XZ7
UXPP8CiFQDy/Rosd2ZWwnaHlyOEleOX8Zfzhd56QrDqQyUiRRquKqyDjO3gkqJAt/36gy1k6z9Jy
8Q+daWG8MKLwHZ88j1xLl4n4CLWbu2n4pbMu4OI2GbZHQFIPW65rKKBZvIpsG8uq8atHVJKe29t+
FKx7uZf0i3/I0DgrvnTZP+Xl183vlGJkZDTyYFSu5vXh8yuxoC6HtI+7ZNQ/Im2HSPyUk0jIAMhS
XDFRoCtl4nnmVQfH0Fg1bK4k+8mPx1PxyXpMmgrSW80bCLyrTTEPJCRgkfYomDsrm+YQGGDRbDKG
vDs3GBoKhfe8z+az49jc1c3nA7/r6L2FhWdAFEjbsekRNf3jMEHcDGiTNvrYt9NJEK2e8rUzQLb2
AQ/3OccAv51RX89NOuGJP4q7sUEVbZeA5FQ93kQVtCmER9yY3OCmh9wlzEvtlt+q94twtZzITB0e
T6gIFJWWbwrTLtcgCnzLCujqH0sQ2r2NY3efS4N6oiOLhYNMGVhvWTskk8jzG71ccEGnd8Wag4OW
ZJF3GX8FBW8C7h57B6YfqHb4nmZYaN9BY2aIisOreDQyYr5Xnx2jku2pYJZyAQQQX1UTa0+4oHEH
quFBenCwWZJP8c8x2BVfWeXAtnyHJXO3mliCK4NsgtrMk2x9tijHRUgmwCMK50G2lSkMJqC1IM8B
UiP/9/UPNv6IC6PmLW3TN8/elpVR1DbMJHd7CmqAX/dPuGq7MYbcBcIYoHP5X0TKS9OUIgY5YWSv
FtoJDkgQ0ZphtXtVnaVkdnqVJ1D7mwYF7HTBUL4evlMgDyt+4LWNtpzxLuC5py88gUu+cVivd0DO
T62i1MIGj2YPKKCFNNde21ZC00W6uLvzwXCDXek5qy9JOXidYvcBn0wZl66eTcZWapqs85/HBamu
06anz6NP9xwHQMBeM/oEpaN2V/CTl68ptEO/QmEvAs58uP3elRoUT02Xbl5KQAbhw/5GqtNJkab+
8fEPhNB2CdoEAGWWXXtPm+HgO/MQx8+rvHHcqi08rqrUm4m015GY8n6oFJa5kJWHuYRaLuJKD8w0
+PjxOjIsufJTe8xLtht7asPKa6xCYR9CbRs5kIXO4HWubgKTptS27KntptgEtmmsWQuzzM3GiPsc
5zjf8FP77voyJguqyt8TuBm1diw3xFm9C+3UdnqhsfypWxkI3zHG2JgDRYJ3ikOTYiZj3OxM7Sgp
S90QlrCUulNZdVK/0e4tRiK3wxW1itELE0gDU/HT14zUcomkSMt4fcxgJc+Sq37Pp+UXILoMPmSv
kTBXoxba7t2eBqiVTiNDAJq6YivjJXZy44gjR/B8vnNbEUpfdhaL7+vkJqUW9RsE3s7nCyKYld2u
ICh9Ln9bByESxJym2DSDe2gM7cgnZVm/0p3Zz0jWaVCK7HGo1kzeoFuF0g9euGTTqMZ6s7VqMv22
+46FS7JTB77ZaMF+5PUb468zuVOMHDunYMx0PvWPST4ljgTAd4CLhdex9l91T0BTZLJlRcDZiX7m
6PFf1e9LQnRUYecZdQHrppGVsaKD1GCSLL5WrqzcNVSH7A5xvWOM0RErE5p0cennac3hGmOY8fpu
nQroxUfeyNqfeMUCWCqtPAN7AvyGfLKqAvoNSUs/Skf43BqRcbeiWm04wsIu7DfXHcuHRpQTpbRZ
66Sly3RP2d1i1P+XSqLkGBXzSccNcTsKf0Z/+PN7y0W7pCKXguYoQhwk7lwfFTrZlxLN9aeUkD5q
CptgJkO6qCbgmVjsl+cGy9dHP63tr1aseelDBZ5zwA1F2TrnsP2f+hcliG9W98VBe0xa5lS6VWHx
x8xqxhqz3Lj93i5nG76eCQtOberujNPXyQ7mjLUoKyW46bLwS0ac23kQ0vMUTHLDiKlXbGQLjazJ
CltId2hfuRhCxY9yN60oBeiCKb2XMGchXh4Cq+p0R0iKOzo6u1iKFFMnO3EtxHly/ZnDhDiQ8OGH
zFUMV0TrHzrIDPzls5oNO3NUbTinToRm81k7rvMjc3WCrKzmFANsifxfcly/VTq5lTZp7ZzZCVRE
rdbeTcbj5kFJu7WCP599oLF3zxmZW0szr+NzDdxe8HhMpaDnIUS/OTl6qcAXh3yj8IiTZlxxKpth
aHNvc8vroo9ZOD3Jr4E9tfzxK9s94da+0YTKSofmAE24fcXIWX7dGB1nVknZvywxoTNgDuF60nQP
ZPXhjzM/zr7Hv/eMqSKjOp8QJb02EbHldnyn5h7eFh4Y8ZBGXCS5N7pyZg+7TD5KJIKvn5Gpm/hj
qsbr0Fm5lvcUh6H10k4svcyibaYyulPwy9GY3AlPqtKLI650gqTXPhGTRFrBTqAKv38V4b/IYJ/m
SS2vKjBpR6YZqHiM8pkR+U98C3spZ85Ar8wtLmPJ9LQTsiCiyG3JwOKZAC6vfUfYvS0xaH/TI1ZD
ocNdV4QjpTWldvkSVmg51XnSLU37wU/7Wwf1wZpggy77rJror3z5YZ988QV7JUYe7xEiG5ZbJMFt
2wiaxQnl/4eZkC2oW7S4bwUoYQCxawoj99V92xyUzk4xv/94M9f71NdvY1jNrCn2Qs8iZ+QmUpel
u6u1UGYP3WdZk+VkMRpmswV5QAPkunQR2MqaBg/Vsp5dW67QdNL2DivNjF3QcznaEIY8t9ZBpNZ5
cGsDxp4m//guNJQD2Eqs25vb8seleRFtLRBSUKA/Er5/0gy3MKKljqMxoGe25NnszDmLVnM+fTdE
yro340BJqOomlAiNUjK7OHzuOaAh2mP75gsCkMRDRGAHvs0LbRg4W7fLu/XFXnjd8JQVD45RjFWP
bkJBoKQpiO1/iw40CNHilUsa0fiJdPbcdDe1xpkysiBFBev6Q6ycblfvf2S8agLxpK/yJDxiChbs
IfhD2LqFbg5X8hqVwhrHq8EwHMkRFRkS1zKfuQu4zNKxdClhKHFI1nYcXmtr4ff/qBx2agMUyVI8
H/AFJ+mvTtnXLE7u/wnv+tne+sVy8/28JvprS3YZoa+29yWqhyuJ8XNdWIBxgpvLVziVUk0dkmKe
BrxROzpuOp7155OVWn886RN7QlG+nMCRet8ZXiNYwnZrntylvJbkGuTvOP9jw6GumtmfUkcQEJud
lYSkfysfLgrJ+9R1pBAEJVPagKZqMFaMjHNnX0y1sr1f3BASlJbcVhMQPMv+iVEnR0w6GV5WAd3q
D6qWaGcWvF8tPRYyet17zmtHwsLUh+Pm4qVI8BJW7dlV0Gu9fOB+VklNp47VH12uiJ71jF35d0tJ
JQH3ZyTg0QmL7yyoIIWWCWF4MH8Qs+10ojeh+ty3avacwsRt+bvLdwPab+vBDksigxT1SsUpDqnv
x6fPJBcCjJFvM+bX4d/slG+f4adbqaiehBwc6yX+VeroqtuIafRvCIgr9QvWhFPTiGk2cD2/ZO31
JuUs9+GsaoXxoF2V/jrT2yfNf0Ty8h487Hucs+FNgVc95MmNuu7yNk3c4MSAqsPzMoe6gLs/WmIP
Z8zSVfW77e2vvsCHpK4dyjRhcaaYYtLPEjAZIZHc0rtA6gutdYl34rJcO5OKKWBTFX7KMUXeH/NM
nSwC7Rq5SgeyWEQ5qkbN8nQI8h7xZldG+GoQ5/X4zy2J2sOvmrwgBzVS51da21SF99JLcnnYbKTL
/tl3VH2Rlx4DPLBYnYX49+SGCgmtzNnAqLucPmi+c28lGfgZo/N2ZN5BOEQSbkZzAomK+Fa781al
9sZwqUx6/ZEi0tlkXxYRFW1F182R89bGQNgJgF3i6eYu0mhn+L2iqobj7zmbnCx5lB1dMk5fPqVN
UwqMSIQSBIPrnw5Y56Q7+Ca7L5kFZRV1fQY913C5s2A/KlckarGDOhZwnIxor4YfcwWbYzYG/hWZ
4NxSETbDFpFx+YqwkEEWy72obXUt91xMH1/BB8OYe4z9LPgBE7lzjFgwN7L5GtZOnO1PEkbMgjFt
U3AMUlF91RTdzlzg6oTzFeeB6sOB/lLcWLTeRWMOilNoJerKbv1IAldBmjCm+UA43t6U8iMAkiEw
EYPNEMvQZ3fFE1ZeXKKTJXSc/3/ZJitd0QvINidozKh+VOww1kb+vG8JuyWG2IMkhGfr1iBlnkQz
yBidxKwOJx5Qi/3doHuDwUQCiFZnqswflSr0EnBjKUHzqCwgHX5fgIBTuyuW+X57JHTi4TCusLvN
/whaynlahoj/4s11EBNDTJlJFHKmR2GcI/LrQe+xyKDmn3TZ5eSA2WWQboPrD5I6ufu4oQGLcTEG
Dncv3deY99GsSgQarngOUHYPW8GvNgm7CzXUr3x4eR6ZlHDRQ0zXPBLzmcvgN6RSpo9JWV8RBLxf
HkMlzNyoXX7jqGCQ/CfOtxKFHiE6JoE3M3eSe5L1CYRndSQu7I3KnWnNLN0qy/fTE0p+g8MsxaO3
xUFOVzd+gIIWxL2OaG8v6/wsMcsiV8YOVKugYGr5mlDdG/bwL4svAih79zq0WbXGGPfF1E2AWMkn
vviFBbS5iV3yFxvFZL28UE53VDn6rvioHqMxeFi+JxeGkwkATvQLgZP8AYMbufmYjURy8eEDbqD0
2k0+mWu04AWrAd4PR8uHUpsqkXEGWBuf949+T2+MT/IZds8+JYYiq2Vy3dRAO2A/h5RGfLNGN6eO
UOyyxMPlaYhhWOSomyVfk3wV/9uuet2sQruC1lZBwNJV2k3S6YwAhsjxWZHGTLLeRcMRhlHnDFl/
iylGVbsOJ1OTcZ4qAE5gBnfq5lmqbxx9W4YeeqYjUoj63+FmtBO9LYAbTu6qm1dNiMKcnnLmu8N2
kT8vv0dz+69EJ7OSnwtRHwLARSp/rayXMbpshGwxRmonJ+OI/BKSuAkdKmv2NHF8D9mHZ56BzSF+
mBU9hH5Y12wbXTNmzlLWyBu2GUp+ym5fM3W/2g+OrCUtlvL8bLmmNyM3L8krHpYNqc16dp8Y6QPm
Sl802NLbJpA2IR+j8T2KqFJLIbZdlu414q2FlmP/4lJl9Gpv6I1Zy4/9J9tsDtoWEYQyuM4rh+Bi
kS2mXBEemcil7BwwsFiC0AIiaAZ7vT3Y5FN1XhGMf0+jIvZ0Vf5YL0JLRpNdlSaHwew+tJw0IjaP
SI/31KO/hYLusx0uv61UfSVXar0zOMxGAjuIZYTB8Le0zr/MZdvZn4F3H/YTzJv+zvhA6uTPWb1z
tBPgO7qKir/gf9q43R1812OgS8etAhPkYjANrtf1bWa8E6mGy5ziRyi2dw6To8F9b/5cpOyp3dFX
uhTzqZQT35qk5GN5AiBC2qbAAkKlbd5gCXLLezYXvPAPNJW0RhaSW4gS6XiLYqX/EZAqYTqv3gkX
kadWwsguBe97O0GVfdlS8uRa5aZYXoindhkeZgPx3+bAMmFRkZZVPlwsbBQIXCNKpNzEwWgXljjc
/JVQrBx9qhLvR54ufjm1H1jrA45PucozqbtCNVn1+2GNgIWVkzd55xN3NegPRqcK69bTVBQ6GfDD
JurF16bM4Q1SRL2SaOW2WwgZ7+IRdVqTPK9XkFWIUk2n3V8ostClzqpppEtHf6Ot65vff/KIGGdg
U5yxdidM09PrtWZKl4m0md5D/LSsOAvscUIsnF3lJd9bNKV8m1w2EHBgI/BYfQ3Xo956epnAYHBX
Wq79pUpF1a+fh0U/W7VVhhXGn5ARJwMHSZ1/Mb2AuQF0OfhNU7qQRP3it+cQhDF/wVMoX+T+fO1O
4jXN14slu6VO6gFYb3klqpk2pW7L9oaekiwbHuOFNa+RkI5VZLw0Ihyhyg9WMY92mwTdL+mIwyI4
+vxPkjT0T/3iy0URFFChpi9t/Xeaa9Up2hYWH4NdKeTKaeOxGS+hcWIUfJ9SAqrNbhhkMfl6dVMR
31EivUs5NJBpF9C+Rr2OYuxpi7gwqsAmrEauYJR8R3hOodPBkxKY6OSmwbDtzkHJrMqcTwMYqXY1
UZub4L0IkgtHf7wrT0pfbFcs7lC6N2wugkxMDyuothH5VqdiSDGVnMj2N+6QVEpXGLJtX6VDYqZq
GVWb9lWtDF024m8hbj3iOCbr/IRSRasYmIWgpsOalSvJMN9KBP9LFdTbqhokcNAc7m24eZoiZpPD
WA49gSwofCLYhJZWfSo8vpHV73rONpKvRitt12qujkGTGItBRZXbKxmk7lrljlG6qUivAmGeot6r
xP6kNc9T1ugr6ZP8DddkcidUI81Thv3vzOTCXTjJg5QhQIEKX0sJ8rrDMgNOMqtwMxmsIAM6AFVb
zHlgJtf8ynu89Cqc6f/tUBfQdkKX90+7jGfPOABYNElKiHSKZYygbxbdnyYtUN0lkyqRF7ppJnHh
tiWEpBZML2N12tunVqt+VtqtzalisS/+Svxg1uNu/s0p0AalissaKCViXWVun6eU3L/KQBWWULl2
uJ7XlR32jR3eep/PVtdF2UX33aadN9IZ68O4sl7lkT6jYltBTxjtc7jfNKQ23OHtylAuT3tWi8e8
uFtOMfL+ECKAamwSI4kGAIC7bwxRpSlG7tUkODIJWP9FYKRDYiwaWvDjKaYHO7nq32MAxOOperVy
aF+Lp1eRhZkOqDDUVVCNRYrKGsYcE+p8+KjvFCXzhNDCO4MpXVFd/7k1m5BdQrLD9WtxgxM4i9Qr
Ni4T94dB2zqfNccLRVYbWpe/zdXuC1Rmd/GTm2iq1i02gQeuzgO2nGFfoy1SViEszLPeaVg5Udqz
afug1chn1u9EB7PWcmVLXvDYTF+3TBwbinh4LH825WbP04XccLf2EXYIWh9q/GqROYXank3uJDZZ
6Cc6TSEwwzZ++Yx5TXrmIJ9Xtl8GqJ4g2DzRVbRDGqAVXgUbDscsyM5SdrjP8iFUJFGO86tkB3sK
7XgVQk7XpDY8d61gPm03I3oocYNLRu39ZpXjpEcT9OpTKL9R890eqqt7DptaqonReXJXuLozWE38
4JquT56IFxkuWRBGBHoNc0amj8ECf9WpSHU+YJy7Cb4WdIiN31qmfdHr+qhmSfo0R/0snBkXPpKo
oecWhI137cd9Id3OKqa7f9l9vW0hoz+8DqCsVCdFLjowanalz5IxTBXSer0sow1t4SMIRCL01TnK
l7rHSN1oQ8Xp1P8ITbc7sC+I+ZHlpZ12zC9WXm2s55+ZGQWyd9bYpci356CIH/SLWJebwMzhPBJM
ckbedx/s2wDjl53/lMsXWp06y3CsQMmv6Jcq6/rC0T87s5mWgWC87bLP70eKzskQloL5nfyYa07F
R5NrX9UlJ+FiP28sMosLTvRTCBvqAA1RBIJe2uuhas2RBZ3mkZDEwyAT0fhKAtcYjbOuUQdd6tx7
TCF40G2AE94sXjhZQAPGFyg91xEqFlqgXeCrtLKrkwm8joEe3MlFhjoAzzc4Wter0b9/SsmKi8dO
V3m0HiSk7hZd6Xoqv+Puo6xOyPE1LQnwgaD6BPVqQWiJ9J9TRc6BhH72Z42Rvhxna0r6vnjDObLP
d4Wc39TtpJLD+z/mMF/2ESz0M3crfCW3cG3ptb49gw7XSDCfEm/mH9YEWmIzFjtVYRcTJf7dwEau
nwgXCoq7pmu+DvSi/WHqzI23e3RtSgSCqC6RDxH0HxhZz1KF8MG09x5hrIjdj6jw55w71so4RPca
W5x8S1o7CXpMFmbgqV7IrHGxyAnQXg2VRw7q7YkzmZeW65INLouXEvATk2UiuPYlw426WCXxdZW8
wq+wOxwkrIVIu1hvoQvAgRpnScje0A+BkRK45FT4HtzMU7Uz4T7KJxIEQqI+EZ5L5qCAHNyYfPRI
zuUlvtep0Bgmm4GbWdV2/1ijFJEla0ai0mFVw/MJ7oXuPzHBoZHwwnIacrGD54NHy0OflXEGnkFu
jX96j4JslvAJ1Dddf8dBVyUwfPawR8nwmlLr9h/2u/C5paAAO70P+5dj+BlNgoyhfsijRe4xcoDd
uyEIpiYVw076EC05RnQQ8MQo4l3QBW1R6f/Asc8JJSikzaCZKT9Td8IdhDUZaF9uR/iBb3KN531F
vEzbi7W6arn/1jqT/3DMJHOr6f9uKcHOy0wfam9sldnOaqhCeNQAVVDvVnU74YHwC9vbfmVZ8HJR
HPhsuUE8tMNHPq0AFbvBumsoE+wFGt4N8IEk5baJrjqsBxwPxg95CDmsR+aF9zg3+vp+vKsWlBTb
h5j8kBwmHPTNDUDuAAK2V0wTmEusED3lBvVlHQ38qlGLK8F3f3W5t2d3Tmk6KO3VVq6j7HUtH2O8
MvLslOfYvWB+nMNeL5W6/HXvXtlBMcMt+KSEXbt3reQrvZkvAtm+0VbzbswlyZAm+GSgq/iI72s+
GVcWvEwIf9iWgL/yZKXr35MS+9Fxkfe31Fd21xwZQgx1Ga9717whFBsLSTbRwZJfLwecolTuKeYc
VhIa2mgjH8d0uqHCsPThHIixlaBu1HslhJrgMmevIwjSM3aIPlrmo+7GK1vJ5IErbvUSfHPkaVl1
YPo1kKSNPlLem0yAZ03uf5N8Iw2KLnf3Oms+u1MGd3kDgvl2eiDWClm18aJz/0uszIUbhQP1BW5z
Q9bV9jFpgNgq48rLs2KwGVVqzDVCK9uDN542YX4+waeGrOIusNVXzsNCSL3HEnD1oTH7IILkG9we
jrGNnfY5i0U5byuF4c0QXrN22BLn2dm4ybW9k6A9LyB8pusAV2y8bv+D9qy4gN/0ohgZff0BeYn/
sZoDsT8THGrFrVcHoMqjh2mEVbsVQ3LLqR6KgFt+3bnlpSJCKOUKwKWmDP7UwHxHvR02naInVzer
HiSOVvYuzBOFBH+XeL8lKSnDIENu87vzqnbjbwkJwISgRrX9TkmrtGNZGTRPzi4a6e5qCVMltWgW
OXEmriz9VBlw/tYT23b1uQufBZSWKJjJ3STyM1qk980I6DL1zh0wpIlh98r8xLhEzYC5qwm3Ql9n
dArCfryCA08qX4eWQcWWfTk5FY9mXAZyvKW2ZBAYwIpTH5CCg/tXcTInM9a+mBfX2i853V9kx3Md
3tZ7qbHil0hO/Kze9zXumOGQvEkrxpqKdhShW8ZKfI71hqGNyqbLd8/pmcT3Z33z/cNkBtw4U7YP
mNZ6P4862P0Hk5TxtZS4LcIVmlNg5V4oRMWRXhaAVWkgYAANd6HLK4r4fajBwzwRhJUBSLiCLXXC
/oHXJTr0Mdd9knFtNKBRERZRoz4742cdc4drZrjm9aixkjKJ3HU1I8rPAPX33/nm79pcdAVSppYV
p+PmTeLcqKwyt0GW2ok6lPljWHOBETaIZArF78GYIakSK5VTZ8AA2bjY6lqZOJNldZi9r1MOWz3x
5pDq2i8fHbVHSN4f08i7kJ7wOTxyoRFN7tXASbbwXpfSEJW0T4UaSpkNAPs6ClFrewwlwDFuq+ZE
NqRN/IhEe4j5PuO1cGDD1U+opSHna3Zi8lwoC1o28lPIgHjL89WHgpInOnXdvWg+idMW9aqyZl0T
JFSSywHDT4iie4LDS4hpMVZxOPvHlrHclC3bwcjbUXz68mlYc3aI5lvhdim8KlzpkZ6L5pqRte+q
jlqIMCr7JqFDBrGJkCevENYWXGA2gUiteRdKp2FYtM6H/Z1mXFyLU2G8ogHwXvXBUI6HpzJSzsJ/
oCjtLhlSZUBv4CMId0MXtgalmdgHQnefNOL0EUDhqsxrqAll3BUrME+OmuZtVezq01DJ+mosw3+u
7P+yqAtTNTth06ipFvoz4XMCN7JfaRYB9e+sm6YMlVMB4potNsbl5bIkzN4dNPMRlmhRqDDL1cJR
Oud7JLCVoNpFl9xD5Uh2wS5AufheGcqZ34oO4WuVWxK/CaeTGq4amyuqa8fjs+KtENp0QSLp9Wag
uGIgCyKuzkColymRZXRNKIxyqFmQzVFcNkvsVLSufRcNSbWkLI7+3UCX+TlyNQ4aGen3TMeCF/hk
FqcLuE9cFr2NgIpBptKUvNV8Bz76O6XoDWWSPYsP7dWsmjU0+U9UMD3Nu+4xQLciF+yDHKh3OIzK
MIQ5J7o3y0IKJq+EThhtYhWBRJwkY8O9SRMnpodRh/gOXiNFIi9Wyij++ewHIgvLGs/kD66oE1PG
vIggP9pbVl0CX+4xTo/fp/R4yedIslg7GbeKpJZn1z+2Ooi5Nc++SIifeFd57QZkiLApHrz9JOfl
noD+6Gdn20n+jaroa9qVrwoyZpRrJh8/3cRYHVGqa3EXKUTjAGJWST8j+xpTsL0fxTOY1uQlcdMg
pGZN3+zxuwQ1WN1qINAMohhvl21APlGOWZEGE1duijXQvNBWKmBhO/qXnxmWxf0ciMhMkHKoQKKK
HFbbOVCItqbhKn3snc0bw7lM6qHlefsT/+V5sWW+NyJr8PdT+hoONLo+pIx76YeLhfp/ehlGl8/Z
1UJpWANM1ZcdX1IAVtPx78QIgf01jVDdQnqghuy+zIvZUo6QZL25IHUTcNCtODBseJh8ZBvwxuBG
NaBgWudBE3hRrV1W+qiKt41nWiOjDeGou9GHMwZoQlR60UagQy5g0u5Eo5PpwS0LNOOZl+umwOZ3
l1cvau4+11SitfOPDZDW9r+Qp59tf7QzD3fsHEsYPtNX+mht4KpBIrZR21SF7jplxnwKBlgxgQyN
ETy76nFXDEbKw7O1UGULJNfSZoEY20yj+JvLLajYfm4donvF7KLtAFE2LDQHLSP2TP0YkR3MYYqs
c4WhsVMMetdFmj385Z1+eoHQKBshQOyGcPwIOhpIzWdEzs0IRw0Vm0ScbQl15440lGgWLGzAJacZ
jqHqWiBBDvAAsjQmSyQ39DPDzEeundgQvlfWB0BQH/3k1tDncz7ACGgNy5UQbFjv3kOsBK4yD2py
3voyA4aM/vDsE5VnObsFFlQErkF32VU6CA2PD9gtBUvuRV8HPPklYQApuhB31liiUCNQEj3NW6EX
GK6A9MNtWiS/cDPTVbXJ4K7q3Qj8OxFbn1v1iEA6XiTW/LabRnsxkaCqE15rpHEt3Z39JApqaUQZ
ybV7CelQJ7fhPuR3cP9dYTteMdV3R8rLG34uwqf/8XFlBOtd8TD9rIliprpe/JjgWr8aZG7K+NBa
hgJx160XUnGqrCwmL/R04j36fVM1TGgvBZ0NBO32XKu7LsE+Z4WLUoaRNhAqwdm3hlGZLDHtqfZ8
9Euxe1x4wnADY3z7doEIpv+ASMxtzao4kHFXnCvDIA2+hNbakczoc46CuaS0MeoOPRc0HYC8bJH+
zVmryhOUWQ86XtPt7R4kbDq6bOpqymFqUix5OXNE5ch3w2KF3EucI5hDhWEP+A5DedegsnSlmmrN
YZ6TYjzjBriL5sfmBrSaMvBHxQVQScYt5t3xFmuCxt7AU5ocrywJJLAPsdKqkl0WYxw/AhmIaEkl
PSGjLsIf3A8SmpsjocmzcM0bdhF6RhTTfuOq9ipPhO08bGi2fXAkT6bGLEAe/elvNQ7MNmR09XNP
OtnYfUr35Qgh0JXXRIzQNKmeujr+g6URsDc1LAs3lMsB79N3wWwJ9/EgdFPkXlQhijenhcs5dy7E
06T/P5ooiAdFvDe2bmwT0CE/qN+aRZIcC1RC7kzMzI7uN8tnK7Kin7BIjWHOgYiIdkIxixINV6MC
g86crQF2rwjnDvw8XMpHfp+IwM0SImhFavJ2S8DG4e5xt82YecvrMI/vKCP7JnGvrP0Mm2+k9Txr
4ah5PB4q5q8rXd5paCxD2Xu6rBWDINlmjbeJyStBJOJpfzAL1N7aLYwFhtYfwm795Atijftm4Lck
fNJ4vbTiRLhWXsbeE2k7b/VfyhqEZysyYOWjXKApQ5MdO9OeIrluPWcZmx0FkSQekqngh0Rut+Y/
mCpPe0EZIDjqP6RBiYqmSNiWCB+zqS84Cy69nOkUTsCJMfx6OXFKdZYNlp2fB+f2HlBQHC6Ss1Ln
I/k9/KB4joL3aLBGvS9PZXV0iEDmiUAI4Bf5nODsFNjD44Hc5grstVAGUw2tnTgHM2QCPrLqb5Ar
GKvYlKPb6/aWpV/uqPNgjpqStSbHQUMcvQpXRl7XW3rzs9iyHLyJVZIaQrByJC2Qn2EsDBCPhbOI
DYnEUFAssdKJupSF23RqNtr88jrG/te/UP+zcEZXugfWav7M3keLA5YirO/xM8tPRHRQCJfJkvwp
AdElJaV9xQsY3ry1xCXSBifMbLGQVrkefwMvgewGxKvpMe2fpUnhcP2z7nD+rcjV4hoOj7yzw69f
Sz8CAeveb39vApIhqDcHcdLn55O7rN+iRPdZN/vYSw97nIK/64A8sQkWTHnlngNYj5IVhhmzc33K
cOElFw6kgoY8sZZ8dmG6GbSLY0TEY4MGWPFuLM52hfJvV0L/GH3BYwwsxS4YgpnQQM7PPsA4J8rk
80HvjADFllm9pPFrOwuv+IeggIyq/CRKoN2OprP1xLI1MY+PE9sO++YSABc7mWLHHS6fO4OnH9g7
BzbolAqDHx4qrNw/YfKHmJ3EwD2h0TArQ0EUIZi/KLaORZfk8Df2i6Ia4lYm3HlRr8qd1I9RpwlO
zKGHTjLydnV33kc6+GfxcPRedZoumzUmkErrKX9wkuLCLUzk8OlAxH9l6NC1/OpW6+SYh5CUYu7O
uSQkd593iKdwWalFMVFHigjPg4HKn4TLJ+OkUNsfGcQJ3JPOk0bl45T8YOc9wZSGVLev1eBZ6or/
bgaZFVkV/Dti9xDtM63NlUiW6HJuY6LYfzWjtK2V5AYO5wYS478iXUqS7GBd3GWQ1ygr42An6BOI
/lbo629pPPfL7oOnaajW0PauMUL52YsReDp9D6WpDTldzaNfElEq4mHFFm9tRVCXXV8+AjCIn1Cr
CaUyCDjTRl5JRMp/07ONJsLpGnRzaZzOsNaJ0O1mq1dfbd9SR5De1ymAcK4yiKGFBYEk2XN71JtU
LMB89nf1PlSLcqu5w2wwPhGH8hJLrm6QmTLvxSZrgVmdje+4m7q+xOCylpiNUsp6aFt9veEkzy/+
L3gNXUUGZbwNgqlF/w3UdawG4+mS8zZ9QXbjYvKUtIvPsOI+SbaIqAFQeN3XOkUWNMJKgn+TN17p
hSp2CvtYf9kShhLCPprKKVt2TW6kLTcrHCHIV3lpdcDYjXjhdMjOhkRbLPUZUdDAtMZp8Divf9Lx
1JfgT+zo6frYxdWLD+H3hqw7/hslHBcGf/kb3epPq6LsYsJo9zJJn0wq7haLuYuo5czKSHkr8L/K
3tb41oSPBJWIQsNMzCXQQjKcK5jDMe9FGndfZbgpD2Nk7fjh+bwAX2q1WdFwvPBRGmoTTUtK2rp4
zTbJWTXbIROZIACn5N71AyommMyCr+Bczq7REImlFbXeZKbgobuB4mKhV5E6n9JK5Q2Yw9dxV6kr
91fk/5pnV91c1c+MBmO3U7bKBjt22BhLFa96fA/M2fFG7/p7rhvRWZu8DA6fs920UzGgbS15OgwA
pVDb+rOD686cViHGanjH9F7MnSh2qPdUfFQYXjgAQgfg1RFY93Q2GgjmRoM4Xblv57Ek2r+UIKup
N99ayRrUBQH1qju0miLme7DUQ9m8Npivr/GzAyU3GQrNbhgQ+L3N0ERyM0qbGHCnlxC/7F0+v1U7
XDC4ES3iLxDkfW3YzYK59fFfJSi2OX60gHBqqLajSCC8bOuHgd5auOjELshpttaodLFbD9xkBPFe
g4+bBJcG7ddzBKE2YFOaG3lQYVEIhV3cBr1JJH8LTLJ9sBnFVV5EFaIgIVo25g6fdZLqXdK27aQU
awMpJOZDRG4B7WNtWZnNadg4nrrrJGieDn5iCyR2aDougL348PT51G4fBx1WCHaQHq4BCjoOcxS3
ecbQu39S6RRWG1VwoKCaOv4Jo7jc7LSPNo4kWAUnBBq6EQVi4XyGdo3BByYRMwi61NiquIPgduTq
/IJ+sJe3Cn2IwjphEj3kDVq3gvwzneEYCjZHJb6hr+ag2ksAtVwmq9ELmTnQsqOwriGKub5WfCkq
d/E9BeGV7Heu2TkXZCO6sqjwjW5ezcpxBNJYNj9KA1ckwzotr7fPSENAJjba+xn/JdJ+td2F8O+s
rkpO4Irk/Tok+x/pVRPLDnQ1Ivgxf2azvB5O/nhhCRX0uj4xXECjkOrGxA24BmEC25TcqlQB8RX9
H22zY/GNIf2b8YQC5qIL0qn145Cvek4++IJQxVPzSn68FACNLZsV2kUvSJMYgY/1ObwhvlpTRZyQ
tJlxb4SXKLXaWwGgghp4N588D260+TtcT2Cr1l47HJpFYLatmi7tRpvi+5Y7PEs99rJida14Rylo
XFn54G6Gm5owk1/kreD16E+aBmIppMJjy9NW1NVdtpS/DlM6PZhDSS7bu7I6L0PGSjCYyUUe2SX/
k8RnW3cZF/NyIE+aYT4+79ApYIycSjfPlf4oxaXfwGYSuOyLUk5oUziqomZpLDk9PDNgkHilDIGV
WqndUyqV8l98Zu2cyi5iXB2b28BLUHffxBshRvttdXuP/lce0kVyVLTSEGfJXDxoKKr9bhaNqhg6
4ElgJUAQznZffouxIboiohw0ZzlRVnvAjst8+1Wci+/HsPbbARm6H7adi3QIlACFcWcOfa45Q8BD
LgqjWSOQdK0f2AXn6BZVML9JJG2bnMON317NHlFI6xlZ5Vk4BojFgAEtmb4wj84KtUCHPPPeO4et
Q4VI+7okgFmtB/LgteZ46QNe8EbW3y61uAN17RIBw6HqTKGEv81qHLisLEZsN9C9iEBT0n49GpX5
5U2n8ab3Cxbjq2IncTZx213MVahlIcMZSlAcj2h3YSBq+HgrchtbB7nHiaiVcdZmgZrE10L6D+6R
GWc0mzUq87TP6gWhtrZIsPyNlELJQsRU2m4qHu3PaFypLxKbGYbDkZEb8Jr9yxNfFMtG288zqPLU
LOU8OE1pYbz9PmrrLJD3IQXH1WOK3B5JvwzM0d2o6O5fa0RZycT9e6HXM5J9DrhuvqEvnx13Zg1d
bX3fcIV9F47rOluPo+LaQ+bPsdglmhIhgLaifO8B26qDu1q0MEwzY/1X3ByUA8zBZtHhngO7MqFK
WMgJyq3snKN5POYumWnnF14iYElVPQERvqIBNZatNk/Sjt+oDU+FeJ+5+6uiQh9kogec6RKpmVL/
SNMlvhP9rGVoIvUt4izP81kDaJTFusL1eMJjjsiSs1vT1RmbSo94Vaes6PT0KuTBfI8CPVkGvdGT
ohMMKNjWVBD8TL4WFv1qiYC3X5UTw1SW+vrV9YiAS6Xxad3zpsBa6PyU23rOE/wELp3YXdsaB6Wc
YuPaNc/r+BTZWzx6C/2DvBJ4KllFdxayuUQo3xZpoMWrQRYj2RC9be2WmyO+WctxaZf0dP3wU86y
6qdtI4WZYq/+VFPDvOFTdHGfHbg8vhAXDuM7ZNDy9jYqaYmJMYmAy9WltmM62qw9uAUdnELPfAaF
PENHHWjJ2rA4UNsSkV6XjaiETUKpO0J102RkZuDwfKaUhO1NQa1s5f0fDk6CF7YwMuXOWK4QTkAB
e3i4/+JT7TMu1z1gLlKQpGmZLniRPqspPJt6baivbAsSx12TskLJtDtm1eaJ/zSGGyC+zvzqV52U
mvn+KwBsgbAkIxjzCOFZAaJtgalGDK8jOQf1M5n6YZv0Y4zwpB5jsh/dMgyeOxaKkJKz1xYaANng
gu8BDrjSQNCEhivyKcNxyNQG4LiML0uqzNUQl5khkYCtXe9afiGMS+p0udMoCWY9lwoRwHMcoOHK
1Om0k48j15SRvmypgqVXH7mrD9Of1gSXPjqZEcTPXT0R/l8kbnH6dEQJI77yQ4+K8FAKU7x9ZK8K
gNOl3t1TX3R1JcszDHkJWaH2dkY8HGSVixgbvISIdpPnW3LsYYAGIU2cWjMFqVNE+yQ4UrRLAqos
ygLBdekxYlJOVALUssjVDako6m2jff5/u3tjcIXWPXnO47Z5TnVyC0VYJol+hi8F1JHqvdpk2y1q
heqq6jCvtU0wh2TgCuT9wU2IACmsuhN9US4qVk9ivkaZh7l6GUQEsnm/9fXSAwAT6kuNFCovlH6g
C862xoX+PpPBaJMasA52/jd3Epfg5ytUQNRYeiLeKHlQP99gwc2nO0aepl0Ne6EydkhOIb5ufOqO
kdxc6knoCG4Sqk7XhEHYUiOjJpPeQkUXmmHLVhDG+AKRGTYkQ1IiTvrippS5RfxHzDNuGacZZzvA
6xeQLKUZdxu000BJlV55b4GoB2NrZ4ZBb9CTbkSz5M7Ce0gK6crCtGrcK0oEm1bDNUtqzYiGRGZU
XeO1scUs/7wjWt43iIYZSsYZpcE7Vmk1CZDd9Tz+DbHSSQYNC+DXspleMFz/AEldaNPd80/hDkQw
VLdkQKYgMj0eDKaFbDlk4eyd7o9WDTwNPceIZ3EwDaHS01akr9wg8aPdmyg+mQdJwTdz+nxQjrsp
EZo2ewlduhr9CEOCZmZZKXB1PYLE2PM9LytT9llTk6NWAB6umWoW9HBHv+F3a9aU2uQuhNSXSpkI
6mmmoAcrask/Pbrr9kY0P2PjXg7YM3Wl5xIVV7EqP+1maPplFRTj97i+4mLfRZDIv18vVlvn3WGn
FoxsfcIlFyHBaL53qBwrmH35JM+64W6tugApVaDZJB9d67DD5gCkHYbKT7xDpifZB6w2p9z1hmrq
GoH/bdkZ19Q7BBwXEWZFWqtNISoUCs9vU8dZSCZfd7vOFfSOLfXW8lNvII8EgvL4PHCmXXk6zRj2
22I4oAPaegw6d1jN7DJnLm2rq8qv2n/V4Uh2Q8wxGB0hTePBLoiVf1+6ocsyClXaU7vhIpY3b2RI
KPSJLkBSCWc50sfhetwFCIEXyDWaAxFFNZv5MA2VRZVLTdxpc7SIq4FagYKXXr8RKYJ7CtPTnd/a
o6p1se3rfgDQ6i1SF4256xztyAdFaR2oTYiGhnWjopVUUL0wG23AzmIp5VZTVp4mMpiwJV42qptP
v4gRlWP4cObqExiKhwZePk05rD6Kq/ytXGXLigMYJNyg+5Ll3EM2wyaIcEBjmjKMv6klM3Jxi5SF
GKCvPWdvF5VXJz4tanr2cwy1kh/L2b9lIC1UHrOIuaBZRr6z0kn7eSjTm5q0IOzxh7a6O8hrdeDs
eu7j70GlSCw6QyeAIlRJSi2Vn3wUWyUDIMjxqqCZbP2WOSRZ2+qkrh0dZy6ba3LmOGf4H5mj1q1C
q/a9yEZzsYF/QoxCjayRFQxgEO2BsWpXs3InpL4k9eow3tS3uDhA9bUtyJURjN7I64RcBMywi1FQ
/sUm63z7nSEC7FTnsClbC1xid8BJJCihG3eWFKvj9fBX2cps2J12WgOnu/KuPAEzxL8MoG5m3OZX
D1G6LJz+SSlRQd5/xy+OJ9ll3qKRpcWodSmjqGINtfktdzP+n3NPSZaJr6CY/G5/6k3Tstiul1tB
VCUYBSpnI9MviKoEtju0siHnyJ/GkeRoYUameqSedH0n9tKTTczFw+MrZYQK182fn2lI1zgyyaHS
p2OgFKi81pnnAvt4/GKTQ+oUNOhC8U3gTKJS9aWrXP172lKdP4xG1hddqS9S86jfeL2Kh1oumJ79
gEr8bZvtjxqh+d8Yrnwy8o6WWX90AWyNQ4g2nWkiKYN7NRFnBZKiJK4FSjDogjkMR8XOm1oCTVPu
qkeTL7auZ22cAzRY/G/Q6SlLdHEBJvzJQkXEf2nyVzBiTMlatjRNPSi+J+b+VyCmAxeXgJ0j/NJU
VCKvm63u3466Y2h6DNCtccmHVmnDF3sN1iG1UjpdffoWdYgZ33Cf8SPqzCPjUjHqEJflzRkwmfzA
uwZ1T55qdG81DXGAcfxvC5ZwKbNSDQvsEfye389hLvrmgpEUkYCWyX8hWw+uMY2AqADNKlxMm5Fc
J5/mGxrw3qYe6kdJ9sb/QzvX+MVdQvJqHWy0cVz5Cf9Mczm2FJdJol4p7KoluWGQz55hvDiV0bZW
hBmbRrz7FnaqxgXKHmN2/P+og9t+MgshDG4Myd+Me/c/NJLmgw+Iy1KoN6Zs93CIIRULcDz3FS4F
E+E/YS5kMRWPRNNlxO+rRQ6ftJ5n3mosnmABbNn2q4viejembzR0miVwAYlkCnOdVy3EsFqadH8Y
S+DclL5zpfsDO190ks2rfEb21IWD+FTnVmqO9e1pK7S7bzPcUpwvvu2UzcFU8J3CLfGoNvYFRScS
A/6BqEArIICaU4G5A+LM2+GZCg6B3vSGSif0SLWYGsepB88oAMpX/9XEHg4f2C7yhW+0s/4yRR/Y
vyBLgR2Fa/AI3tCy/OFOuSrmkwfPpVRwmNJ9S9As67de8eaVDgl6K3Gfsu88wOZgmjWTxezchnpG
SwTPRSiAG5GLjjJcYA45rk4gK7So/oPIqyL6rWc/iDNSLylCiR1PqMotmIpYhjo7mGqD7iEcqd2J
CsJiU9lTeQh2Yc3zz2S/Phx6PsJiUbPWlgxGo5hjzIuWGnAtk8cnjJWHYsO8zwW7btjKfqTWr2SL
LPegHaGSRAS5a3N/7YPTtmrKgXa4grhDmwVENyuOUVXq060yAW9NV0AY5wagg6qF36WpHkyVCb9b
cf4X45eRNheGtQxttbnpWfoCgdpHQ8l09nlow/p1ZJCe+ylQhnwqoXDq8sITAK/gxOu0dlQlanq/
CWB4R80vjEPzj0SKe3yN/d+6TDanZSuzW93gLk7fKNJ+gvnklicBbzolZTrT0s7wrrjCUrYEXgBD
Xh+XaaxvX9E0tFrtifDuToaFEFBxQdIP7HLiN9SlSiWeLKIYiWR9FQ6m8z8fuM2VX008FZxENPLJ
tznYaeDTb51k4RZ4YKkAlrKQgYQGwIL7srXLeDKrU+cNKemf0akogUZXsjgxGhtT+hAY0dlx4rFV
d5pujeY9pZpcRyo9ji6fjOjiUHJp2fnRr+QOVuou6Gmx5E2R+Tl2TNj/jXnOERlvL4HoIia7td50
mTqj1DT9chnneGM5qRJy/tG3kt6HLeUs082evZAC8hXzCcWsKL+dKZD0ZD9lVyf9mZdd4tayThb4
1uv4U0+noIHIJQ9Pm+I3EEzr6jeNWEkODT/oP/n80PSnS9c58jbAPXRacpomLKXtlnFlvpATj9c9
UGguo40vLE+NBfVtTt77/fl/xETEt/jbvjtJ9Yp7SlPMRxnlIxm9M2XwNWXZo+qTAjHv6Iq46dIE
21BanrgxNGMbrWc1Q8OQoMbfRZk1JS7R9nGwYXlQvUofnFb668yUlSjFggNYJ3CV2xh8huin+p4W
NbgxY9+R7x3pE2vP4ZjEqqvPNEgXcDD46QoC2EObapGELwenPwATTWCxoEJmOpS//UB+02QgpUMm
fQotrzJcDL8QuYgaqX4CbD79xH5bhTV9oVxx2CwyQrv1x3OEIQnIgxCyT0t7QEiVIsEz/stuR+4h
/Y2KpqnODhZ+vrduG0gkvrrCh00+NYYjlsUvRs46dITDXnhdV5oPcO5BKlpNsHVTi0dCa3104GLR
TlHxEIJ9aIqZyArwEqtUoME2BsdSWoYuvOY0SxmrFJ4turH4Ba2l3HrvjfD3gRO/ZSQKq32WwwBq
KqwkNWFqV3BrXswzNekss4YigMLkWBKxFxB/Hfe5jkAlr+1E19BKeZwMd+i6GtRrFK2qgaJK9kNt
WDQ2gRw/IwF7Y4lJ/HptqiDHr2oXf0eXa0GrRF3biLcE9XKQXkYCCiNXxBjoB6jWMrELOOQVp0OT
7uU0qbx83uxglzeSj8ygW5Pz/XcSVYp2oI4PfAbeVQ5TYWdJ0rkkyKjp7z2EF8SKfy3lBwiwe6J8
wXLb59fDayA6iTyAjRARvo/gHjTKEIORVh+qYW9W3aF7MiCZNQFwDnwSnf1M442sM5BCGD04BGkD
uqFOIqHqH60MdMXpgTN3mWYCszEfcZXp0Lm7xX/P/iDducrXzjkJd1Y8LaLSp0Iu7j8FjQEwBzYO
vw0+n969r7g8AB9aI6Ur+kDFrxxVFij5C+lTIZe1DVCD5pLnmkwBsPeam2wAfJNO78WCODtY8p7y
rBq7KKd37m6YCAaJIBUGPlRkLrYMAM4B4W7gNDNDtU4NFYKozTtNOEg9f2RJzK1thtfH5o7VsR/t
clsFP/ES3BbrG2PrEv06Ug95C1GBDNOnIYCxIuX3/Ya8Rs3ddQaYr/LJSh/ar19TOaQi7dNz2Pmv
d92+usss1XZI3YNdp4ZQ7AJf9CT6/fikBHyCsKX3A/uPERRNZsWveJU2NQNw/H5NFVBLu2e56apy
UferVrsKFBHdatYfNHWfaIp2Sw/yT+cSc6uZ/KA+RUhK0O9ZivIzR5EMwJNPWBlamDRk/H5QO//e
A8T4vDMW2qaFMNRsmtMu3ZmOiPRb4nc7/aMsL4dupuyzQ8yfhvFYj6RbXYa9/p2fGohMMhFaUHat
WNx5QJv9hWmykW0uL8t+CKoc1CvHJJGAKNfeER/Tp/XVi1ntD+wlG+iNFqLbUDci3ALJWJFi+2+T
rU8GJxKA35uPYYVETKisjugdeNIpOUnQhecC2BrxXfJyMKGYpLanKIe1+cW2sfFOdDmoptlIE5d/
jpVl4m8ScmSm8Yda+5BjooE2Lo6fJc8N7A0oAVYDU0L0ISbNGqnA9tLZ0SHbTeJmT8Xrk6RU9F0/
Rmx3ReFDB3jn0dXBVcAaSMYs0yBf7REKNoU2/iWs10fl2nfgOlzreGON3dz/GKbn0aI3grUV3Y92
hzy0ekswpyY8Uy1HhaYyZIFjHdMH1+u9fIgxYkvLRQPIVXHc6UKoXsNpJR/371ZYfpuADeRZTYLs
EoaCT5paJtfYKp/ys/6zNk585+MC4TEwfAHi9Y1p/tEoxsxuM2INnmjUdchqc+FQxIm60DRRDaxO
skUWvwHjonM0h4s/5PEoxg+Y0zPLYLLJkhyX1RnvcAi8fFWpqkDBbDcyPho31GMXIQxDppeXAjs3
bJq0q9BSG9apzeyCwXgJXenmDa+Lr6eUrXHYqEtfid4LTpyVBGJaNlwg0u+ovDOs90DIVXO8ixPz
p/c+oQyEdCsqL6gGTFve2PjMeYoC93FFY2lIRPntyTYl/OMxe/M8uzhLZrM+J+8dCzE/0xKAljRu
mv1ydpyCoICNFNtcIBLT4n3ryJH1LllLDY3kIlXUSSAmb57w4i+CZLZHp+CgqzAwHKqaYAHDFbHJ
GkA5b00yIY+JyNQTaaz0gEd9sUzRSf58KYBqQvobIlCammDixKzn0/00LmBe/NLtDKAh9j8+MEpA
M+EIEXKfxaWMDb9K1x9yFBF14PQVbLMLWzaIDPiO7DZHtOn6o4hOYrMA2/LPkm2zipCNYrU9zSxe
tOKek3L2ajY5MK0EWyX8XgL8wG7c/+/gWg4Dvr6VHdM/luoV4o0/QHpDSjAVBZHqd47GtlCFE1i5
6x/xb/BbiaEs3mvw/3VWrZhIst8ietc88srXiO4NRoPYOCNcaC3JGvNKuPpPruhSK9Li/rxoTFb7
emANr1IhFqrYOck9010dKVyPbjmfT3Rk383BwVR7dm+Xx5/ejB5oe0XH1kVyBAjPj+oSsRXIC1Un
4N0WnrI5nikFiRnmUJ6ViQJm0kINJKb2bPbBy1C3OW3K4gyS59COfEosLfbG1Qz0IaJ2hupK5hXs
o2RBEM8bHGOtw2vMYPn6t+FDYbZShYpun5raV9bXGP8dWyyWW18efilscinzznXbRhLlQ3HhgKZ2
lWp6W28sbjz0s6wFUvxd6hBgEm126fOyEz/PNa7Y23WS0kXjlAmK1DYDyYaVjt4nHA/v7FUTYsID
KluXcJINwy4N/DT/wukN6tNLeWDC4BY95YDGdUSP2do2usz430d1Oo/iI6qOfAHJceE5gnQco3Ld
LsBf8iiPJo5YzKYWZLhZMcZzLzIIbwG1JIatlXg16tAHy66IvC6YPe4YlMiuu6V7uTI7zakbtDD9
dOxzpkEGiucKwAYrDoYA/WCD9vorePrm5g/Q1azHWGxVdFycnNiZix6tGg9p5SvteiXzd4Goh9nP
qujYdkGyfPB2MmitEN5UYM8zy+acAZTOv56/rzAWmqtwrOw//zq9p/e9mS/vZww7U5KGcOWQyIK+
yzoBxoQj7RfFOVHUV0732XcwAiTqHXLX5SBtZpTe43IjI69g0LucLIbbhqg5Y1E/pY8y2kDKSuif
Lw9YZn5pr3UwnrDOW/2eU450hF463pANjE89tpa81w0uP6o3UIEs8KghD63cRIH2MHEfKbZVHPe3
xN4x3KGErGen8kizjIXpJPIZD2kXJYi2e0Fg/Iq/YhPmfAeUU6kpnbP6Pi1+Oy1oeOflEQ74/rJ/
X5Nrm5FN56T2w1oRyxA2w5CNW8neJqTbXeN20WrzYZmzlXRrPxano06i5VsjMM8xVM/1YC37yxl/
NI7qjMj/Ltpu1g2RDK6lquoaah+vN2CY14OyFu99aoIdqkfi/gK53hFnY/aS684by9bXoJ0X1q7i
vjRXj4isqzyb5fIj/7nE9qNEecWXgroqHRUQz9xnvlo9qUVMZddRTPCh2N0A4Xk6D6BjHdlwb7Sh
dizNopBT0x5rdzkry6mxWWzHGN3JfrDPA0UVGF/sM9o6dR3ri2iIJlj9TvBCxr1iwg0Tgstc93BJ
FvGWcSJXqvAosEC8eipZlMxnXaK7E6eTDweXY+vf458CoDsojjowoillVnBzhd2PwXhXNBqBand9
g4XhgxkcyOLvk2GckPduG3JGXO0SuBlHj2SA3RLeT1dvCCOgaYthnyjRQFF4EnU6Y5q5LrmjoaSl
SE1JGcYg4Zy05GkqckSosY0rERbRU9gRSUJz/simG2IQTgfXZFfl4ppmiKFd8KxLC76UVwTn6O/0
vTjGGAmK8v9MEBnuk/bgWU8DelVwUyIyQagp0D0AiL/Km2PdPJCX1bk4TLmPR6OfZSC/p3y/jxiQ
qBdiEddjCkHXEUEfVj1ZUd+FuT1chWqIeUOzdBl93ecXZXcrwF6SnzV4zhr6kgeoYyZ6qD8XI0/3
JcOmQGlEHUPkFxBFtDycFAl6YjIL/MincO2tRxQeWx9H3/RmDgbsS8nNXYc/uP/jpUkkEsNsl0A7
K+I5V7RxovLUpdIpXC6Cx31jvzQHSV97AWezmkgbpPVhfy3pa+T06rOWGBG0itr2PBr5KcGeBeQg
CkqI4NkBocWsnbrMWl1ZJrNF0S33Nq09YcjPbgVc9+3bVXUc2Oe3JsEi4RbqsEJFDSkTN+nVqfzg
F81IEuQASV6iKMmWMt3ynwfLpyz1SHgzl0JQuoGUsS9rxq2LIGMd76rY1ZUwfmYzDFDDIY+wigwH
VioOakZ6ZBTXfMyxGZ5OpBUp2MYQHXeqB8l9LHLULA2qHo7v+yWBL/j6gKZvybo4czFJT7rQ1Cky
SngD537oPbnEKCgdPT0utRnOLGiasazRIqNkkYhpElYyA0Z1/H4y10BpKeERFr44zZBSyMju5RrQ
/2wqfhfysBUZmfsalp+iMGS7Pxg9GUZ+hu0Jngl2OrKD0jJWj12RfP/X9eUvjTPlBowKkJg4VdEF
SuvAmMqCQmcxTCNf/WQQH9OhFG1iRonx6g+8yZRPaDub5dqXX8EZxTD6Wdjq/ikTHkIEMo7+uyBq
81zgqEw+cX5DBLKln40qN8uMbORF1GDl0oawk+32T3kTkoseQw57JiKcv502sfQHrG1kTRkjYOHE
wfwrM4PYov19Esh7z0ihqxtDMYTT/QJqBGrQ0ywBqLGv6Y0oPRLgAaOnB1suU+E7WXJFAmpIJojr
XVmsqMdqAdTZO2vW4H0w2aFzLBXC84wj5BjcK36LTghZeew6Sr6W7WtLapy/R/h7qInyUBiVsaOp
E6P3ZXg0JHXKr8ekF/x8fbuEn5bMvwKZZBvDC7YXOctSa5aCElzmTocuq06Qu6V/JCzGd7UmEODX
DgbQZhjni6kV/nL4QvngwW13kNf/K5Bpp4M9VIBKiQJ5kiDEeAhjCMjzUGfB2w5KEXJUYr6/BYpF
AcMYuNov8tNp+oIwR9HPE55qL4INACzTM++zm9x4bodjewCsHOXMpD9lqtSqHbaTRmp/IIrop4EG
uIoCR9+v/xSQCNoIaBmPHtYqhryHTvKVFUkbZaYv7UQ4WXqd445jD7Wy9M6orEBGoN8wQugVYRQw
kEWlMDmMnXRcQwOMUgmuzldW06a6e3Xrtl8Gr4opr87tmGh/s6/nuM4FPV1rkM+7XjDMpTUR5kF1
CQnLi0ASBD1QQHvklcmc5H2Sic3O4nltYknLXVuV9+7ELJq1zE+Ed98s6BnuYNp64eUeCF9f/ym1
Q68yOV5glz6nNZsMSd42AEC7GIasLR9Z4JRcfOih4VhKYYJH6nbbZK4kEbATZwwPbXH5H1c2a5Wq
liaUYpEl9cvhZP5rs+KCTROb13HXfrVudOFHdey7GfIWeukxLn+gNM10Mux5a8tQa2GzQtTrGEzX
VqqELjRhFzTU939Ed2DMDxz9WdUlI6P6Syma+WMkwcMatqfGr1YU6hdo5iD5X60ZKwe/hOA++zTB
BC4giDa18NFVOW1aHMtuUx6d1pSgwAInemVHpyJxNR83ESFcFebNfPtRbfU3+X/weoy0/czjQr5A
+amIqGoulI4LFaScN1H/cSj9gfPTwdM+IQJR3JjRvuKcoQrfk28+/BYCMwgrTcSgjjSd02UXcL3a
4Y/EECOKJ7Puybjgr9b/JBkH3zrWfOkvHlFZ5EV4X61P/dROS7f92xYpW2Pd5fzVxE9YIWdItzlY
qP6xqxZ3TUzL39Q/Nh0BeUTiJBF/b3/9Smf55YU0tm3ba1Xtd5Fk6MYHLQlaNBUeE7Q0fBvueQQC
46rFVDC0eKN3RrsCcQNqWq4X4LhtxPDATE/0qK4aLZK4G7ot1wo80O/HzFqi4D++oc6Tv3mOdEB4
PYoCpinHrfn9WI304tmNZG/TXqqbzMSVmC9EUcf36Kue/T/nuKqVXKrMh8yPgOsWDSsXDa8W7W9Q
JiAMpAq3HPepEj3EoVC3TBHyTPOUUuHNYpBfh9jqSz0+1qgZPf1lPWdeWYDjCY5T5XTkTf5P5X8a
hxsag/YUdLuQo6GMNNXst1oQ6ertZpbTNTUQZGewx0KhYgipCNS3QxMEDQddlIQK1ba1ouqCrJPn
7MbEJPqyv37IBlvOKKgTRi3gzXd0P+fycoR0dEy126Nm+Mez/ykgi8unWyonDC3YdvA0DsbqodVb
g8kCTdS3GONAr5JyFlSNQukLK6sRNuRTLivJ0Vf8OvQ3dkfSl0f4TvdDu4TBfgllnT+RezAFSJWS
yobCtCC8YUJd5zBpDo9fVWYOPgLwjqHwbbQ80yhlNa7eKzxO/SL9OqCYyWa4n3VbTuM3CPhnb4lL
23tjOtChOvvacq3JAbbq/eNqm5YHRqjdbyVhb5rRVgZweXFZPaNjTVoMPMaE2rn0djAD1sIfUT+0
L7o4om8oyZeiuW0TpkC+Hcvz9+sZyOaScIAzSqgrovkBgMKdNdgZ+hyLLJJSV1csVzrGbDagyCTr
oxX9QoZLKgYR7f4lUb0jyctDH0KaBeRGPJwfOhMEoq4jkJLRCo8DV1EajXrDxtIib1U5z5cCK7LS
PmQpAYhQESLY1/9ZpwTm7OYJ82Lbi72tP/dQN5AhEQjRuNnlW3ber1n+s90hDBD1vCDGdeMqWlFG
RUYUXJeOziTeNwJm5i6UbGulhqKrdNsLWK4eigEbyCTq0ZeJoz4ecnmXZyIveiOVp8o/KiY1d+Kc
jhIfywiNmZmF4DL2Mdcq+mwgqZ8tzhBo+lXqm0errz+yyg4Qx9f3/QRnPywQbgNWZcaOuIyY+ixp
6m/y0h3DbxDGoE5zEu73+ttYDyui2WGBIjd3NoxUo33n6y9MwhDBZNe7M8nYRXRJFg82i0gyUyxe
p+Uccy3I6Bf4j7MA2NA80VA6SRmWymVgivMID0JfMGuGNrYS/rgXezAFQo7soxGQQ8CwzOf3q8Wl
RUKuLjG9IqI2bEuUXz/G9yUnhiDQwnIyvLm4UKXzpgRo6AnT8XgCksJ7QgdK+UN+s4yYx31FBR0O
Jkd0cYKUH46+zoIFVHdNNu/IW6vNs5CD3+YZFvXtkb0yUc/QpDpCYznRlkq+4npCrIzq5C2nNx2U
gyCJphU+1XBihplnODsnioEe9LEROvRoKm5ubqiRo5V+lDtpcaefBbnZ3HGEPBT+lGyS6YzwSpcr
4eQhQNKg4tqgeNYO1SEvsw/ZPAPoIVNgw68MuKNVsqs0ZaeH2RKOPLwd/F7BlmcjD8KLVsEgnSFb
514YP1nYXgd5g1fnpN5oVFZEXn32rr9xVTbQJ9giMGJspFzbag+cjQWZ0cfQkceatuh8LrdsxFim
Z7T0MFyn7gKWcXeIm55hHe5spFI19z35PBC4o65ldkrcL4B0bZ4PfqaPbCI5ODKMGrMap48jwJu1
GkoF9jIXxD+GFKzTXXb6PQSU8y3VPq/v77qLjOvq0wH8vQUwozNxaO+RrGe2uIDXJEq2Jxum2Rdx
8xStixcUSApsHWGXRK8kJKNnYNQ2sbjXKBPmTHKsGm1THlKcdQipRNkPh8WKF0dPWKXTCAEe3C2c
GQBwDn0/4g9bDrO+MpJcNkVfqVzKTPumleHERPH4kmF4OdlQTNRNJio6U+mYgaQlssWnQzynj6Hx
WvAj7rJ4h0sSUfi8PJoVTUdQbM1eyGMVYkoXqMkggen/f2BWvIS+CaC4BeSVktgPgMY8DEr1Rk1b
wndO3a8t9PG53B4IBadlipkdIyt7dRvHU5plS8XN1qGOAIY6CaPHPp0SLUnsJCCQrQ1ifOige6jO
3i/io9ecoVvlLEEK1kXAm3tYx3sFReT84eL2bkHEqI33rAc8ZvxbSf+Wlr2wGvg7TYS6Hpft326C
xRABpTXX0Z3qtTA3G3jhF9KDcXYlg57/J/XkeFW8GligD3Pzpntvb8/hmDX8LxaYdMUkldXDhLBZ
gepj5mFXCI17/v6NdY9xjHhCYtoksx+CRUTcsz9FlkEfIlDiy9efQrLTfJXe8Ipk1ANpUU2AmiHd
NSyQ+YpSm1shmg0GtUit1dC3tDf9MeI93Kh+ycbo3CYV26hhw70J3nmAMBbIS+Gzjc6UzrvXgnV/
hwUvzirI8D8Hui+xUKZ7owjs2wL6U7kPV2VCIFtorBW2dRi3+s0CAjiBbfjrnGKYrY4e5+Eoekh8
ODo7DtMQhW8XV7Cm5TLYNEOh3LogmPjapSd4sN9hE10hQmXIRAEIInOJE6rpfg3JDCwOAqORE9HZ
tt0KpyehkJXHZPCY/Lzaxi6mXautqoZv31cYf0HwNaG0AkrqQ9tl0Xk6bqsBr3DQoxW1f9DsXIdi
V2yqX8HBHiAtmPGT/K51xCiKgtvBBcIJnqWQuJXliTsgzOMVSEQhnBaWFW2ZIRRg6Sr4DnO3cc64
LANhVFNP3XoU398w3VVmTQgrTOqV2aMSG4hQwICvugol2nBMgUXtozEoftCjuuyFv/F/E8KgG6df
Zz5eykfvi7UYEv5fVHPaeipV1Uzolxn1w8uOyc0ZdyL//aMoZRVA9eNkA5UVTKHvQmxHlZyfN0gh
V9ycyzBSWAdYYGJQ25XnI3s4TX16vOsPK901GtdXR1svMojrStvVY6HPrJi25X8yE3HG1I+YpzP9
FGyCU6/5ECzpQH9rkvbVJwhhpc9n/4BXGRr3K/dGXUbNxw0e4oYsFbAFfJPDsd1xeqAxp+pEXDe8
0siFLuvw1jFohOEzBbSt5FPinbX9tw3k0OROfcmAvBs/YUfSl0pRRPHWAO8dmBNEH7A6xSLsQmcs
BA5T6FAanDcQZdSj+veAkR523kUXivBQDB8I1c3qT3Qdg88VB2XDhUZROnLMXx8l5WOx9RQK20VQ
YUnGk60IZikNWq0WeUboY0APssDm/yLYWLCRP6xsis91JD14nUNcmsxBAf81+gJjcCzr0JuPmalS
lfUJeQzQo+iGoWGHsTPu2bVWZtDMwXcjTInrL7AQakxHBKTl2t4u1w2ygdLosrxeXSrO4bAw9AJU
ppKbQVOwpdKv+l0Bjhz9CMX24YfgXZ2bpH2kRCi1NU3OmwqcSB0JMl9R6t5tLQXEoUxYXpiV5a3m
WUGgEwKt6mB8tC2XKwcanp+cWdS0w/CGEA+UYMEqEqD5ZeiVHAfUhYBzYf20jTcj9jwNfMHFI2Fn
tpwPD9Ja0JFIImAVSWIko7AOZ5+4Vgj8FeUueJw0iD953IogEqu8Zc/uMKPTAa0qYeWzeWrArJLf
q71YjGubl1spS2bMYNu4xHJ8x6/P9zOZaLTwJPOd60zbjaWaxb9fNyiM6o0ley1zGfEeKgYsfxBP
FmGQBkZVBTzFGtAbST8nizjHhxXasd8JNEgNT4bOgl5I6fNZzL9ONQkeK0Gvl6DChkLlWwQ8y2l+
bOv9NXaZeRrNLXqKz5pOmgd78UMAKaEfY9cMZ8muFE+4e4FGuAVfJ5yj+wc8qDG4kr5aD1MmqzhA
WiZaarNcv0NJOw7WhN1nHHg2ps4vbVxLVEw8u0w8R2PaCkEgxWWmSBkc6FYMQXmxQ5QBQJ9C95hN
N8lj0K1WmD9fIGPmOs63wUsboOS4uKbR685+CUisM3A71hLCI0ZCLIBL1PC/8IFwG7g3DKMEPSFu
tQGcJxyicFf90TkO7y4BnpYFUcAGHEj8FK6TwrODy98r+qMlXWl6gZi0AkhWZb76ChEmHDC8wlVF
V1PID8KCEDKs4llhxH+/kp42hrkQYHjJms2YQ3RlhjyT4k4r+b0hTpJRDVHrqjoXpo4q2tt8Vp72
XPqhFhstt9VzvxE2iYsee20dNF7uFvBiBEySOBREj1rUwPgOn4PS2lXh0jGlad6pASFLQ8o59E5J
Qry8nQyvvj9Oup78JQqqYEuFL+uBnIRcWlIUPzgcZwMnDsG+zgz5DO/aQwa97jw3h/jleux/niGi
QxjIuS8a6W6ZW6mmIuuiuFsexcDcn2v24vnGPKAt6BQUpCCuKU8IzC9r60TP0D5PXli5SyQfEzSl
kVDTXQzqxXW1WtAiH5qA4biGitL+pLl8mA6xJrxhBKpxYZd7QVOn7P7ePEALV7Iba0qdUd4gvFSj
fknnD6e11Uj69WoBLPde1T+V+6LKYuz4+QgEhdFwQ8kPrTrVKlGti5rukfkMQPDG8Miafdo6RNAk
fVpYmaXadQzpCeGIr+RFcs0S/lX5f3rvdrvLlIQlXHChP5MKBsfkgRVGwDDGgfj0FZeY0LVGDO0W
9vrhIzInMZVaI7blLsmGLFoqLCOgdmU7JCgtKnHu14/YX/uu6jYJqkRzdXPiwbCIJeuAD/Jcsb3l
n6BQlvMyT0X1MEdyBa0Mu32HQmyoFQGWNc1uqlEkv/2CgPomDzjhZgnA48GgmQz+SZytc7Ut7WYF
feuBTHhwiX9C0MVfMJP6fZItQZtBhbfUTuK5Ok/+fxkyStfIT164HwYayt1wzXzXCNTCV6SUCDtf
FHkH9ArunguaQDa7Cqz6ven50xDmEnDI+sVD5uNBTbDXEDwMrE7x07AwNYpY7vqKKVlh4LVb4U7X
hNtz76Vf0TA8RfJqriYWWXxdyKORJ0CziUFudl9o7Xbf8MKykCR0isLilvEsXbr5K5MDweK4tz8S
rqql8TGo/kj5V2M3bKNnktZ3nxgw+sg+ynkNKGB1fsnIsrXJNjwi7NKXmriX3iDI0a8aMcVPHq5u
rKNyUGheJjYsbko7rwbOlElTV9Mi0mH3Wxo6mHZaOLxTX9tbEW0DOZSyqFH0JpE3WJFYB+vgYURP
iCp5H1UQSwAooFCYN/M/3iSxl240uRMk0KaYHbL74Q6prF0HEyAYSXKtGW9k6jsR1ElT1R5/znVb
rQHH80JW3wDdpthJCLDi05sDUQD9pfZjMWWoJF/mPLYGQAJJ1fSuiUXu4lxzX3doxjPEh4P6KIXl
yWF35gXWV8SpjQli1KzXlAX9/vYu7JqVwaRDOVpO2IpAE/LTioPIy2HAU87Pn9YTl/z4W25Q1/90
DNQBeVNK5apK4ziaKRXe1bQblAcwwzRRpX0HlfOMKr08Dh0PuXnn2CsGPWudhFSKNJ0Ruf1/IIo6
OVOfvkmBhBzMH/mrU6ZH3SVx2Q/tfwTSqACYjDZ7wU17wuFpqUgc9uEJYXgQbxdoDQ/uaAv9mo4D
djNK1DADgTaHiO47i0ie5DbZWLr80TXKRnsh/jx83ulE9H7WT5d/nY3Rdu68LdFDQhegFlqHugu+
tjQGd98/g6TJ0/AwdGIywwB8mvB2+tpiU0Y98vtz5b+tZNcUIYVrTUzkS6/cDN4eH7Cf6XUpUv/V
aMoFuiTqspNIL0Julr4gKvoR07IZI0IiEm9j2dCe1v0lhErAAjTkBmnOXZ1s+h4P9Ln3WKEh8/nA
QnFtvYha/NRQ+v0+Fxm/lbWutLOkNFpxoc8ETky20BL3/bneGUdtPpOzUFlUoOGMZIYkKWAua0hy
P2b4Av/Azt8OLvn1Q3pW8IGkJADFekLydd8ZKQqUrDJo+1N5CKWF03tLBisH0xweYJshtcK9Z0By
u2AnOEFWgA3KGHV4+l8Jrs2jbpV6L4SOcFziwbOAhSsgVBZ4cisOAl3X+b42PROe1gNLGr8XRC4d
np+qSoKZaxREzrW5et6FAo4La0Aic/DY2XNWz/yWNDOECBXTQlbfSCsHk9RiWsRG/gWTgiFof62I
lpkK3rnxp00XQGTBDuwXamyQpmsgULZFT4wDO7FtEISdBe64E3pnF9RBRbaZIMHHNvLokSsmRcTB
PPrJh0+9DjRVfnnDS2AlYoIx8u2TYPyewKuwFtTqVX5jgpf4eViUl7AKxIeg23iOGK9+GxxzTpab
ASdwAdT50TRCIC8Xx9gJ8yXqakYu/gbL7fbDaGu9aFEaWqtAMgrJ4Gc+Q1EPPmSnID8l1Qrdo+a4
Js+x6BRkHwBTbd8+kHpv5pUw09zUy/h3ea/dh4Z4M9B+m6jiLFMZ/S1NA+qGyJv/uS54kxG4uv7t
ZOUfWzHxHfIdvOHUCdmKeUOn9NIUNCWDKZU2HgI+PLKc8tNxlJmEBZtsAQ2jp1tQydNGXul1fqIH
FDwIJOS4eJtY2WKspVgM87VwIEVzPtOfiIi/pPjLqKSHBo2OAWhnOhQlg5ynQ0HPMNDH8uJ6TILS
QTMrG/Dqi164pCn5WVXxcBhoxQcI/NVCslsYvmkFFpgQ/RuoYAELiHsrOeLpItNaWErislIiR8WD
W9KyL4nS611Fg3wMKes/W9c2l5SvseQgizd3zrDvm8xP21B9hhTCHLwdFBvRMIQ0EHHrkDUlF7ls
YeyrKk+kdbq6SNVhi15cqKiaVw4CTTArcIB7l21t2vmfBuxxe0wgczrVUfBJ8PkYQ2oGnXhHytA5
++RZfiAE/plWifbJEufKhnsNs73mghq1LfaID6Lx1xD57++XzZN1q0PubIFATmoaj77CFKZKRazv
XogdwHohVWwNExPbuHax7PGUU335hqGPgsW30QKOxrtBNhTbGsjy2FPl3v63vkuYEIH9575i+4nh
gHYd5JSpBYMS5Yi6+v2vBCv7x5YVP2/evHl35fxuU+jeVraFUqcGSkc2wwkJ61tIaxhPInZFCTdp
GIvF+rPPiMSRrnB7pAJKahTUdniXQYJhriRZUvOvkU0QiGf7Sn4QZ3KkEcmH/oQBHhFqFh5aF+MK
QzoPJ2pwDXWrIp92N25UMrxYuN8fNrI/Intpz5UC/3zgmd+k1l2bD7txAgdPMBq4SrhGRfkJn/yy
b1iMyql1Nd9jGSigBIyM6yqrRiVxFt4WC3qUW22dWj6lXlx1K6Acj88WEnacxLaKFIpBrjxA1zGW
TErgPopOoUZOWcFPVPqibkgLxunDsDD7qVRr9DbVqblat9uLSgJH/D1E1d8nBV1TCKV+8Hdf0IBR
nuzCLjcclxV0Y7TllWX208mAEao/2/KwYPJ/dSsqQobn+17WtFkq0GddMu3pHWgployr8sluV9WM
xJTYuX9CGHNnl+Mr/eHW3kvNUtXMAu26F8bcbZ7Km9l4Nu/jKOAC3zs/DPzOa50JGFIYIMkKhwjc
Wqv8WeTWdHx08phbPibQod7NXXMC4CukOJnctuSdTh6xEHHji5BYKez9NdW+tgU4nCo8LapsN2oS
T8n3H6DXoxoUpAuO+KaNMIVR1dlU3pdcId/u4jOs8kmRwX7pHTYlbRpfAcvmb3IP/sNIF1VZuRPc
GnY8dt7TbcQ8iE7wmawQVpyFATL3H58DXJmp2vL8EtuKyjNiNFK1+UfjYSeZPw79t+dUhDAOhITp
SPxk1gYmVgu5KBg/40javxBtS2XtPRhYMsmjnXxchFmMkQdn4s480IJNl+aKOnMR0qgwIWaycgzZ
3tf74iquarIUi/VHqOnD1TlVq89yPX/QKqaYH7qrMkjtVRmoRLcSFAYPD4+PThgB159UD9JI+udz
RtvOisGjhn2FymmRdPb7TKH4qVnEg+ir5zUAon2Mqgtsicnpwt5XLLX/YrTcp7WgRYmy6Pct6P8j
dZ++2QvOk41cy16uQWkVKNfi1DtOFnxuDxS/shNJomAXxTJqaGlm7SjBiF0RDA8bwhrlNmmwnaiB
6nqQ0Ej6g5GYrp4VJQJIbauicQt8Jef+HINqgyDcsRIU3X3slW4XUKT/0ywz+mz382AYX52IzrlD
X4MirQjvM/hjWZEeJ+sWZijggGiAeAFYqeStkrImaiVGcmvWBMnDDKO6TM8N4EnLNmCfxIjd3YD+
ZuB0FgEZXpfnte9eqR6t9cKihjOPJqIwGKNnxx4GnrEG/z4rFHrRlgxbj6Ll9GaNsMlsNgDdwIDd
LxZ33RF51KT99i3GxlNu/V8O/9y2rQl5GoHTR81lCmN3qW68+f45fa7DrE47aqODtdgAZtsNSJRI
m6lwidAkpwfjeGUzFbO/b3rDnN9zJmZf23eYKImmIqVunQn3wVLj1jPKjn59HhDKUkQXPAzHUi3h
wJfxn8yckt2P2OVQcSsubhM8llVeHghUjz8SNko3k2eXpUxHXIPFRUqzbwBHfADVRTDsqGfHSv/Q
mR5jlg63rMg17Fo+KhcxhA21fM2SI6Pp2LuZlJ72F4GzRWE7FODq7F3qNi9HQHVmcWMt642eLyq9
fp0V4ZTmkBYClka0tnxzJJDu91Vx0Mz2p1YYJr0/KlUjK5nRXqHUunb//XWhXOqw4ouHFdCARKGr
JN5ubH//7XFcfHi4F8sJ2ZMt4ycF1TvznZedpQ30iCeSp2YLlD9gMo/fboiKl2X19esbd8RYxBBl
NQ/ptU60U8cxpOdw5SeFBo5M/xTgqMtXKCPwrOC342aodmbNomZR15AlUesTbM2Z6l9FV+Id2PX+
7+4enlCjR8k9DO7LmvyRVWKl2PyhhLMZ3s7PYhAMQn2+MwuxP0fSRlaNAi0fR3jXMHvOUQ33Jlhk
MFBIkTisofnyuyTTR10OsW+uVLVlV1kAbCuRVfYfauEFckACOhIMvwt8oofXXJriKri45i+NMxYJ
ac0nbLWSju8Nf2SKmKuUfMM6zeDPC8JOAcwLxLum2NhjVoKTCDRwU1DL4FhAUTYfIizcYRYdxuto
1n+irLpwDX5cYLGJV8FP+26gesmWLvuptBEBQyZczf3si2Se+wWNBsNgByl5Kz2Oy/hR1R9PA6bF
a4tzrJ2nUcsvb0m+KWA//Si5aB9OHWJHDsK/2Bu2PHH7tghvcRISQALMqxsBkvDQf4CTReZGjzx0
LqIDhLbY1UyQzJaFcawbgSKsj2hPpBzz7lVCSoW5tgcpLhUt4cKgiPHsLN1Gj8czxMBkSMfHQFne
/EVGx6IBSjs3BnNUcxd/fNiThNl/HVQyLhTID+auPDt7AkEwPTXtn7AK8DOYKNxZx04eZHwTm46+
/dmAro+kC54SKYO2T0jevVxv3KB2/82Z8/CB3V4A7S5Hmrr17gIXLNVpEmc7/wEyxpoQ8cn1Vbj8
B7k1f6qppPiNejOT9qtZXyg/Is9RgR0aVRsXxAbguV75GfBel/lsBypye7jnMth2mFFoQoEo/FGg
MSFUEALLf9+XPYiXz6XfXAIwceDVVsb5lWriSDcvgqROor+wh7LH2BySgo3gN4oK/yrRIA6WaSAp
NQRC2D9DUE5Ga5dmXIPgi/9aQXIjK9xCl7+8YqQiOEWQLeNkEywQ614xmU5jocbp82GIfWwsfpPi
R88DP+7dICvJTwdR+3rwFLIiqYStbTXKyS+3DCrdJvuLaDu6MsvfJLtlhW0yQ9Zu4VqUpTAVlUBn
/OK89oIPJDmpwwM+aXkCWDGQsEnuKDSYWq+n4zL3C5ZE2CmlkuYxrt5lpUWLrTIfgYFSC82GdRgn
tR7C0UwmO5eFKAKrtxuIP02Exe2anT0kE9ibGFs0bfgLj5WzZq0Z3r+LT83WGO+KwP01tClBgqVy
3o7y/R0aO+6hT74C4IZwHpwdVXRk7noT2+z3r7sWnbiAHfv/3pF663L5WZ/f9E2He4LWImuXFO5c
yNgkJhZ8HxoodJAC5jMtu/NNJnLEgjhp6f+9t8Mh4PdYP5Np8F+bjCUTOYk9EiiGn95wZi9VZWDS
VSD0FLPD2IsTZ4nEdpjP+BIQ/S74anoqE9jpLYKOgOrCs1kOJddNs8bddXfKKdToh7q/Jd/XGxC/
93Y6EvjhSli81inW/mYBuih6BmHZZtYj15d1BjyzSPk4kxuwlBufL3asH5zJc+JtoZfXMne/8fXy
orDvJ54pDfgqPwIR8sKTxRre3dWa3HItVVac87SvIF95npjcZNB3m6ndieFS5KvP+Uel5eZ/F/WA
8O3wEwzS2i+3UFFh6JFEOtMj3hlhwfFzJsMyyRnooImcjSBNsWqbRAl1e2UK0soj0YBCcYw0U2su
FNqQ8a+1ou36Y5mryj6hq+QGZY3bIvgxqnqRNWNyYo2kkqHFIMseYwF4RtSZfKtXrvoBLv9h7YgS
cq40QZnbrWx6dFrnzUaVDwpt/9ROlHAm9Bjh7WVV6KjzQpDkkhJUWQ2L38Puo7DzpZQ3S28E8Bx2
rF+0/hqR5bTIev4NTRnwCuETq0KxbMvKApgf7goG8M48w+pmMCsM81PybBvanZBgMiqMjswrE20g
0ykwIJXg/4cbVKnzb3H/gqK/5LaozKNv/h9yGiVr5xOyXIFvAb1t3H0XYh3e8EYdNIEIHCtyv+/A
MQ2/zMHBybNXmDFq3InkQkVYsVO0sGYis/hWwtpARy2r1eVvmpNjuXLjVRyiSd8nC74FOGE20XxD
QBRFKvtyx9zWEmLebgXV5Ym1B5knUf7XbRaB32rSp3iYNuW2x01hOKj3A8iBPt9ySffwRzZHrL2z
fJr11b4zUz0DsiTO6rOlaJtb2Vuzcpdb9gCNRSBHhI3AucHSJUVmCEfrQv/XmL6DvsOGxCrbDkWO
CuXLGw8Um42tWKitX5QlDL1AhQMNWmJsLdZU14d7Vi4TUTJQV0AtBxm+i5X83aes7uu0N7G323jX
NspPttMZ3SdM/VRFUoeiCKpzVkM00RPUzdjBsmLsn0JzgB9nuMSYioY3OI8bSpLG6NMX5Urtj1Vh
2sh1Sk7mjXEo387b/wwQ3fzGROyeBBhGbgS9rDCnn3ygKfn/v1oQQibEofBoPHjjNy0zaxDKJDDb
sD/z2o8vQqMmm2AracRQ/LBFsOjqv5/dz+uK9HfWCKaBMMSdfwGeqw3bD5dpT3P96o1vWIvrDwuX
IlrhPSMj+Eyg3OlGW410NhsUAF6ItVcgHhD508ed2j7yu8Ivd2SZiJL0ab1YHzE1pSpjzKwLjwKL
k4MOhMrDy1VYDnS/Dbym1GnoE2D6kmEKQf3iMPLvxQe+XQoJtD9lQ69b+ShHmgHx3ZT+gajP0ptx
mkca7ce2+Ce4NzFlYGDRueJ5xhFLcXB+pvbjcbqktMUlm1vtBKBny3XTkPZibHEzykKfcy4DmBn7
70OFC3m0r/wDNsxLcZ2LowtcwHZ5Vqsq6aUb4iE6HyGg4SG2W9/0x+2VLuS4G5MNp4yy96un4+BC
11ncnDxTV7au/n9+Fiz9DaClk/MIA794j05ln0OBpjhLO7DYrrqnBq+9oOUwy6qFUqISILSd+vZY
/cE3ARXUi37dHWl/MD1BvLT5DAVqHiF6SJKOIN3MVVRSqaF++oYENcnEItOOdY7ya5or5ACW+qKq
wnB5U96NbwPKwQNXwfzxtFH1dgLCV5ExBwRSifmWFjzSAAbft9040blhtObdfjbtixVyOQWimFub
vnOgsIeWN/UvAtxlR/CsXp27+l7Utu6Qdz4oDACFxeziq/u0mlv8tasKYZ+tbdQ/AgstX7kj3K/i
d+hZRAC7KPYsJ3FnOp9SlG8y9tmwEkpjFceoJYh+JK73uPpBeXD7eiTpbT7dSkt+B0cFZ5tw3YCA
rY/Lv8ySvDC/nCEtTDbQ0iZJxhLFSaA62L+K6ArkgcF8s1tf+zq7HJ9HLHGxNcm5Njzp1+CAaILl
JvM1+OyJpvfEMcbK0Werg/zkqhMv2QLpxG7wKg9r8+n/MyO9TN6MIuzCOp5zRsAhbXHKunzILh6m
3DiC21wxD5Qjr/JbVi73iMTLNJaHgBf8xBb+Wr5xVwMHmTXsU5fH1cepAkCeu3lhUKE+sfg+uyvR
FI77t5ErHvzlROHjHSHmby4HQACfuV88piNs80qwE6iHMkcf0Z5A+LemlbxthA23yx3y5y9JIZ31
NS3oVEW0fbCZhEcj97b6z2eY4lfFBwggrXPQnj4zD2+GYh+FjVRrmRWhOpFOIHbmzzC+cD9SdHG+
1T2SnK88UnSe0owHO+SRwUGEyEL2Hmd4U8wlxDUQuHmMlxDvZLLSuqYlkh+MdA+UVu4OyVOHWzoK
CJ2zC9N6fOfOj+0XupqSsV8n1txvGvYctnzknPRWBsHpz+VYjKvZ/8fN8vs2HuuMjaxDjMjITIJe
zZJit3AkEE76KGCCF+klJ06nWazS+HAZYLocSkJWKWauPoxKPx0QvpX0YbIu92fIxKOEXXmxMtIe
+keitOGUBi4gnePwQmmD6tkf73mJl1SrYtcwWSdD7TVv/dzz+NlfZ9qJk3S+tKjbYCmrvRgQVdEf
j7dvgEBmJou/00KkjP/gE0uokPw/F9ksUTWlYqMhX+Xb4Jx5wpXaUbcQnGrEuycHs5UP61KI9FaJ
aqfPKyVQke8+4vby7pcSzo7DbY0jYLABtlHp/0O3BV6E4TfV06Xz0AlyMRzcjavdRPefAo16OxWA
ghGIzY9iG+SnQJYnKv9eB7OAGngP5F0tDa3GmM+mWbJy67Wy6vgu+LIinprkEmK0nBezlKkBDPC6
Ay+Qf/nWuaaKdCVW7axtVwFEnWxG/MY3WwphP9mz3pvj8X668quodKpGUJxJAu8CONpPrhjoypd5
GpB337BDD+WBsg0Xn9iln35dbW9UKBQ95brbNU8jFVJdvOgoda871IRx2EhzGUckQn0uO/WZpkyj
q8+c0fg301Q6Sr/MWIwOPFqRN3ZYVWM/dXxq1toe1IzgfrFLneXlCIRjj+s9gnvcd2jGC7euUJ/W
XSm6sHNQiylbDuU8cmhXR4ZL3rW2Bi0HpfWV8LMHeo4gsjOyQPZmWNOjeod0I9cHRtcxh3Nejfuy
9fC8+BybkW3lJa1tfX+ReuQdpViPZWT7vu0TOgxltZLNBFVWHzsu8SrdqPoTTzVEn2sLBaLd/2tp
qe453hSQmnDG+7B6EtKLjd17VusXflqv4b+eHI1suE8e2hrkTCj2otVdv2ABBl0r3YW34KQOqYMi
oczF8efF/AOOtR+Y14MFmHgjnVIAeeCYiUIupOXlQDr93y7pywHsHij/+unYk8GCMXT7ls0ffFsC
Pdphy6LycUxOzfWeKX+U7/ZbK1WSAnj0a5kHHLEQqND7ewqTWZjTARNNFY0P5nAzde82kC2blGB5
9bcdFlLD9o/pHvrxvsWY6ZhCOwxucL0XL6rVmuRgGi/qS299L7gwKAu7RRBD4Vd/oXJ4MyrzFfW7
s7DW8HMt/RBhnzMRxUi4jWfP2FXA8nnaUl2dbVenNbea795Jvzf9wvHOmECes3w1hFeGhYgdu2nB
A8wocNefqCyY7aN5csSnj5eyxAXupQei0TSyooA9A4ykVH/8/3F14NyRhsztQiKRbWKIZqCH4G+/
X0j7sRWfz8vRqOQ5YTfnWTpsudqIDDgWzGxtvMkFImuFp7vze7aJOmaXIU6N1drbN76LYv4wYa/v
V8iKkZugXbWXBGnIFmD54Ek/40pFX/RcEIb4LsXAyOVm3e97NsUfIPRhdzTTSHPYWuN6iSXj8FgX
A/Y4JoX4kGZh+lQSLQoN3eLjMCIQrOw6A/KXDO31aZShdBrpg12iXc4TPikAL/Vsk4EHvZPJejMB
y5JoZ/Xum9P0W0KWgoKSlUORYH9hYca4+cPyd5UBOw+VUbPJjYhQHzdVfvT7fsmscn6kNpmZ266a
cux08K278YY9uQhit5b+434qzLzLtxHq4Ss55PT1eTn0+vTKEVtvdF3UDUrbBd16ek/Le6BBd2UC
T79uC5CLh32CBCilxM0o4i0U6COvf4BOgMAyy9wix9RdujVuL7N6PKtNnMoeSaJBjS0pql0pPITw
FU9VP6H1kVOlPl1oQ4X8mnb1oxRf6EasZ8Tw3CiL7ea7Y7rqLOZEUGe9NjpkxCGrennLBzDr2eyq
FQuebW6wJNNX7yL1C8/j/CnksKXbbz1wuAQ4bSIeso/odbl2SFmdATXHsBrk4FeS3Kps4rTnvfm/
zC43RQ2Gm7xBlvw//Wo27fva3knu0+Hkki9g/D3yzXvC68hDkcciUpS04J3+Hw6XWicenoCMD8+q
LSMTo21HNpcTVEBTnccRbPfYlr6LZZCk084kwZaNAQLu8AnM25nPDawaoVyO0JaNXSMXsQDnKkRf
eyJ3KWtUcq4GoEdPMPmjghnrqPd4HXu6q6tMRxn2ze0wtNSmhfYCL9bKIY3A1MCQafcm7+X39WpC
/C3tWmYmyHsQMJJsV9RdbsSVk4mi68Q4p2uDaCQq0CrgvhGbNf0XADDs1glQONs0DINEtByGO9he
7FcBCVONNZ3q5kyiimq0FdXz/cWdjGL6U2z13L+731mT53XhpTV7uwcBPov+BOUZFaC727RyJWgV
b48BdD8qJaE/iStlHp6/ZTTQ/83QpUv3VUsqDfocUR4/O1GOb+pLde6ZFn89kVVet34SP7PZgu7K
fSqKK5F+JivAHxFVr/VpPWV8Ap4PQs3+y1uDTptE1AtIz0dpvGcqfrzGdlVSFYAsIVxqOrWLIapp
Q+XWyy2HKoTR4fVtumjeu33VU8Z1iQoEvXbD3UQX6RF2p57aTM1oTUv/+j7OR1x6yKfzBXGy1KJ0
BYWtbX1BWQZiy4e1dyVu87SZTk7sY3ZFjLCQ/cRDebWigRoG+YpGVa6JbegTqzXXkemL95skxk0U
MoOVFvUoI3eZqEkssfbOMjSjoxU0jjlLD6L3hldoxvfyNMfTLUhx1OHIPxudRO7Hs0RINPyY3bzQ
Z3q4mC4zOjMYKwW3vASliVAF20biHT9cYPEWPpxIC14TFMClOVzlsfzGLIhTlWFkIzr/X37G9mPm
ZHiM3FPHBJjb4DKLqxrVLyWIzdg2iWyQqu8aO2RFrDBPJ4iKrfnVu20VLcx98k50GFPJCFIvX0mz
rnHzXsuSIbPQ9kXop9b8G8Xvw7wahL26nTHKABsL9+HcU+BT3Kn3Ghp4JCmSuHe1BcOySP00HSYq
p2OEPMr+10LHywfszeUG8y+/w1it0XU/M+OQ9sIaRZiJYIslcFknYiva0JtZNuqSfARjJ2Z2WbqQ
8TVtFsi3/toJC6by+poFoF3RIRlrF4UEoS+Pk/A2RREHet5uOkywjsbzvPJyiQd5Fy0dEXfpQYBW
xBq8o9+JtviWV8Fsbvkpmx1nV3xTtWn0IdJSODyYvR/vh9KtB9LlKd1jLJ3/xVdwEu/4k3aAsndX
t/dwU+pl5zN3o7+2M31mEURclC8fLi2SCTMKwD8AgTEId9SBPNkherB963MMoGkFNTCCcaY86n6A
A6yg4oBTyJ/8xL9K6QiaS9ks32hzfu+nTXYOTrK3OXCDuwlWIFJ66rgaDpiy+cz+WY1VSeAZ8pHa
06NjlqUUYZYOWQiSGOJ3pSMaSUbO+9oIO5ZSu2tY+iRZi5jnN5od3VHyMrm245RrJAMTADD/5fhr
MeICrYG8zA97urseI5OaZcoLt46BTKri6QbpZpcINH6WbiY0FIjgcFv+IcgMs2r0tJYo6ytX7X5y
l96Fp0LS63ebOJtQa6DPTFm1Jk6bEIpm/BIPkGR54n4kP7VhaLZGxxceEul67uLEeapgZFyZN3pM
1Np9PRs3hXDmaIWA6bsJL+uX0GqDjYUkKdUbwh9XfUpu1r0mql1/YG6e31KCe9ciIYrCwwjSIZ1C
xZ/vFR3gNFWr1/qsoLmfgvPHgVFvdxCprcw8sz1caMkKXkDPhHHt0BdFtcKuP1yTYMKflhcNiTB/
TfhGmHh2//BOXZR4jb+9RuXmulPpu6m1buZM+Wa3A9Yd7z8/yFhCbLKLFwYXbUQ+iPHTPIRqn3/y
Zrsjr4SHy3PJ5VPSPDVzrjqCY19/22IaNm3z/zb5iOqxId69yYntemR5Z+tkFx0k8rKZvZ6E5nzm
0kJAd6QezbgLBZ3vVxhR81M1aSylWE6d4ZSvQtZ7Wp0yoS9SEXmfMYb0MB3Y8e+SeRffGePyPN8b
6vBvW8efz1Ljtfheb3fQXnmYonD93tkZdKG8n2e7eLy60WvZ5VUeUrB6fXJHRQwUAjgVa7SHhy5T
bjYn2xV9/MNnaWq27sA/cX0/ziwjAzTnFZMtHndYM8T26mDeXTiKwCz1POU2WULh4yeZkCqAvk00
SDdp7Y5jMAV8zjdn8NupPw55zKmCGdqwk0lx5f20KfMH3aR00uA+cw3TDfjCuycgWNYJ6At5ze6j
ehpbsfwFjpbxsLJUCeEuz+j/Sz5TOH2WBW7QNjKFiy+/MQclV+ec2E7yRs41iyAz5lghQTvRWKzv
8Ddsq0ksZqTv+Nh0PDW+7G6z0g4Zw1Xla5DyFF3q+kYXaDOphW6c4ZIXq81rYl79TdVXQIBzZHMI
TwkUuMaTqR+lOb+yJ0tig2YMyFalrpeBAw0JO9E1MDuLAedCqQVG/V3lHvO3ZB/Rb4MFzTutI/hJ
rHF/EfIkrX3dGSN/KFse36wq3cB/ljpCEKD6iuShR/l23wOWEACvuVfM90p5s674qqULrK3Y/Z6k
EqWaesXM/zv7gnhDcPc5hZefWgxzWEEGTZmk6k+t9hnTVK+frBDvh9/q/u9lI2xmW5JomAgeKKbV
zgLOD36riL1l4y8AkoIPXu2JDiDZ2ZTgd1r3Isrdtef+zt6/op8ZyMuyDfyQV2KPjENiHXINs3kq
bRABJoKkQ8l2a7l1uGYkUxHKg3VKTBIHF+coUcqT3QWcdgEgLufBmd5vnJa2pcgcmtyZwf+fy2Z+
Ag3NvCDWb4Y/hmHrGPTpVZpwdy0G3nassYWKpe9YfxD7aprXXI+hUtYE4SZ/ILmf2o75ZDgbPQ0Y
f3yR/DmNI996o8nqF0jaWr/T/S+cVzeSXiJGyT02l6R38SJw673Qr1FE4wUyvIL8csny6tCxNoVV
Sdtvc9CxV1SsRxoBSy0oyfEu3GOp122t981qb5X4VwA6mQnDEbLRyG4VtCOvz6Qj7IJvDH7Z260K
opPpCtJOEZ/cWFv/qsJzWH1BKb6GSs1QAEwibLb6Wtm5NX1HqbHJzgdUaI+a2jYUuaGNdTX+K0pE
LmpAcyFiJYeG48EpRqmoNB65nR9X583U6jZgPpFGUGPv2rQhUCC4mTuEBKI0Qaidi0BwtVqOOp+J
Q8v/ptIiDPpJ4qQ//cT3Vgg0uogfiCHFEon32t/l/kwyBsZKp2zCIDtYYEzmrpFFYfzgEjKMz0jo
zT43wLfdTwn6fUUqzxHL2GeG0F09hWv0mU2qt8nnbWpF9VU67y0i7dg1DP46JdGGZMcol60jPn5R
/JifBc8XtmlYykOViKt35vWd8XAYotXLUyr8AnHi0p6iwgRkWA9joJVRHW5UjJM3xZMk8IpRFO4G
UZY+O9o5mQctfSCL+6LdVKFQ1cK1D+AWb1s/cOFmxtp/OxcluO+IuVU8nIlGta8dt3y5nJOKdnTF
4NVLCXFEH0t9d/JvZyKr1WwYTj7PTgoy3wTlMRZ97eZ7Gzc5jrAP3yPVWjmlX0P93x3oBhsBAZ92
dSETL7z0h2typObF5+gIb++lvSEeQf/d5ejHxzIeIp+Dw5JOXg4LlxD5bDaE2f4zzqZUzP7/IgWV
mgQgVsAGY/BkNO/fDqjWlhQiYwGHqjP4QhRG8U9ac+VkT/FRr3O9P0U/0Ca8Cfcx96BmlYBOiHx1
N58tjjSy4LB2PzZXfwaIXXN9AbPFM01Ckj3skF2aGiEMF6LGG89BUFleE7zMffAeeY2OhKic9upC
l8cg25+dhutRuBtAaZFmQGDoKgxPLYI9WIB4wc3FGmuBYhA4kus9mPd5s0xpyJ9s2U4uaDelx60b
/acCwNsrbPIWoKWDgnKtOBeevu9iKm05eLwa9RplHxLs5qnzvU+sDfmW8k9WmwcDmCIxA6jXgIqL
2hXOoQujl7/okQXz/f5jFWTjBWGBlzSJ5M4zunnh2Qi4uo+DzmImDSToH0khH2+IR/rWpWqSYX05
hjRMfgZQObRLFyx7pKl4ioEl4WZ5jDR+jJaZCNJsSZBOuTuX86VjSz5zg2iSEDKwkGYr2kt/8rTV
WhYK/3Af+IK25QWbWnVTzf4p0DH+PU+m8xLEcb3sycW6nAieypUrXmoWF+t0bn2sb6EgsBG89Ue/
XZSNAt59w2f6fF8jleF/cYgmlmbtFbyWCL/jrr0WnIx7JBb8zh5TIR7hNc6XXN1L6HHKUOOCgU7v
kDmcbnuHv6jNzq8VRKsPjzKN4Kbvc0eHo61UIvF25YZ+JS6GkgE/qG/+x05AzNvQsw44GLjLlRiy
hU6A5h8FnuA8ZOTpxCBXsEFlTcCLHCuUgeblMzAMsSyjMgGzl7grEJdj7DXtPh2DlbM/uoBqTaF3
OE2zr9tR0p+V1izYEN63WpoEInl7+E1ty5GSuq+ZKj4NYrdw3BPGwAF0CATpWJl28rDbxAMwReTh
UNynwNpF/xU0nVrEUloW+ATUOwCPOZJf5ulYIUjAw25VpVBBG1liMv6yAhjk8nwnqUMBM30sZ6Av
vdveQoBM8xBzpHEZ2t7FJavT1t+YBxdSCsTcT+EE3Nim8GUnimrk8mw618KDvB6vBOYOESB+l8y3
7lOwBXGThV6/O9pPMKEtEcYwHV6dG+8MUqMzSlWJ/GthKuRNfLFshzuWk2LR0yxNcMYGV35RVOUZ
ieNqf7O2Jd373ZDlFExIKDk24fAB8Woa1P+ld/CRQlT/mM8dZ1ANy4wpkG9DJbRVO3CH2//IUWaW
2W8JusyGbz9aD1NqTxhhXU09CVcrFztQ7wPJSRguzshyMmaQBcF0b/Fdm5YSb3Y+9GFhENMVDdvQ
MWyPjcByjkn3sV6sCHauihdrev0omxyYaiL5/RZwegW/8vE0tbhfZD+fw8w+ql9a2ttX1a5VINS5
Ss6XQmLHekijeNyx96Er63AUZYmJbbZVgvljjtRLhARkReuHXChHmTckXyVY/mC0kJdqQ1QQGumt
VFSrYd5CmYJ9hGkReBHWY3UoJ7sPjH4w3Yc8cybF+l90ErsC+ujJj+Jf2DHY47lGEnfvO6udX/76
DkiW+0G/jAlq2hoqcweww9u6fJiRZHIW1q3uul9/FCVpeG9la+0D4RfFjTWAxtLcxKLeoeEm6ahQ
FLO7XlMw5a9H965M9OAX50aJFCYUStwZGFePiU28n1k7dKD58XbDGcOTMmGRadz3yyRYK55hpz2o
aDcXEMBFdeNGE+nlJBZFsnlMuMybS/yU3fkN4TNlnbFWEa7gV9o8SL6B9Njrg/pA0FQrpa+CUVfW
mQwfclTIwBflC2NwLdXCsqnkdJ33Vgt7uTwh+s57nciP+6vydO4wCrfDH5M9eCvQMZQYkXv9zp+A
mkKU8lvcA87gkCqVUveTJBnwj4UzSaCoi6OoQkHkokU3ws2fRJuXuBhfEzGkJVaClnMozryVbvzq
ejyna6n929PZSA9Nv2bNihGnZgrqahTxTjsH3fpBAwn9V1gu7/Sq2pdQ5rKIGseutFVuDMSLUnTk
DQch/xE1UFitqSuHEPJejFnWDNWjb2BSUJ9qolhjD0AkLmbTJ/U7LcGxB8y+OalM7nqkxVnhC9tM
+zYvvQWlznHj4QP/jgATS+luqadaElcYyrPjx44fYJzxPoz+CL6kBfRq0CgeltOFjdZL6Ptph40r
/z7OlFE8+AnLShO7vz/ZJOKlu9KXxx5BrDSF3ZeyYGQavBiXykaBeiV7abiFMN2rpYxpp72bpqbp
V37w0dyr/yqDpsqTRyEf3gFwuFNtBj5s0y0lsTQOvCvRUT0z0O31sMG7FpcX6q0i+uFIgeEhHsCV
bcLlPhZvn42ImokXeD9by5MmhfS7mstJ+lyhJsggR/8A3JZrU2bTqlrKSq0a15kVfJdP32mcxH3e
cLQpgvKh09dQ9oKxveAnR5vSOKzc6JTZeZhf+zM6rFMp+cYQCMv/diBnLzCoFmZ253s9PTUGGmVL
Ijl+0+xb/6T9lSp6Shs2IaigGANtk79KQUV3vnyy3K/m+nBd4kY+p7vfMFk37RCoa8MLCBVA1HPg
BTvwlvyofPoz2d5ATi47xpl5HV1YVNvTX3CTt52e+6siLSe6safbq3/Vm7A9a0c/KDwzOiqgKo0B
08KsqBGw7Tnd7reBfpilOzy2pitE6InNo0wIPzHYhK7KHeVdtLn0VeZ2EXcy3xSVwfpg2UdM5m3+
Z0HqW8of+ppNSZTetdPB8TKNPCm3JEpnfd1L5M/aD93YcnZ0BDFj7e61F1V40I8pUFcxXgPnO6B9
OlKE5uKdKQGd6XAgf1bFfq+I39WEEhgaNiH+xMgaHcbWrDR/x7W5scQJimjo/8yww/cb0zIiZNd5
Iwh0krYJV9Vib4lNMpwpnqZXbpdxehRLSpPtXc9RDupFKxr8iU6hxF9hZmLjO4DXvWL6aPT2ZIhg
40B4H04HGPTqN+DfXBlC6orKiKo3UpBwNHjlyDAa3e9Uj3cg0asTpXdMK9ipcjzNbNMw3umpYNEc
zRPy91Hs3seBY3YIccaX9sQxcRqzSQZn76ndjJ1n/T+uyony5kPPMO5qWSGbB5owi+an6UqM5Z2j
T3BTC5zk38IgwaSBueeapQpPVF3pZrxTTYrJTLkpG1fhNpG6kkiTH/A6tj0eL8HR/FCfWGegnDhI
cFV60YEAm8rSFIdgfXaXdnK++ls9oseBZoaTI95C6TF6OoxleKg3HF5L7VzAuXoe+4NthPp2NlmN
ZaWsBI7NuzQYWEfRCJFpPfyiI5Uuham9fQI4+eJ8XKLccU8PUdOXtr4SrXmNIC4Kkuso9pIzzb+Z
Xz32hUo/AdaK5laXrzFn4RfM34xhXVzj9DPMdGE0iqL2p4bU5zz8uqWthL9ugagrM8aM62GXk9fd
l22p41r0EWOFW0xKtN7ja2rMT3+/rkxsKRN/7Sy2Rm9flFCC2ASfjTN/zo9NgxBXkYyE15ON9w5U
6IfyS+T7pfc63/xn2EqkDCj8bT2vsHJpcnxXz+r2/yBBXtfkXyhEgxscc8N6jHxoPxFlZzzkq1L4
NlMPz/Kxm0l8098TFKavcze5of1iGpEhu1KKqqnmpWLQpw1V6ZCAexWH7xAD3Nskqo57sAY3O4qA
wDljQK3ZwMERnsZ1YZ9xR1QP2eiqsjvTXkMXDtjymImXHQ0wTq9nNwfX4h1KkWgkWT23B/3SMrcy
MZUPWiUrtTXkmBibQOA9/N5TDrmxoDaEsjxkvDDotXbWb9/ObVY5PoS6kaPQ7S/wY3XjQ/49qeh4
/L2gOUUvQA9qo0DcYrntVp36EIFHuQ6iktx5p0yWxbjWCREMcdjgq41E7WPotLaXlr07ZhVtHNBs
QrNxflHPdytk7saTUMomSPR7LDxoNUbQaHfSgsam5zM2PSat3WsgsilD7c7H7nqEjiYCkWf/HnCL
zAc4KafN1nnEbYWLQ/JwZA9juOdNwyQeRXB/DFQ+c2/qOslAyHXGgjIw9/5V+aYKYBibXgEkzWrg
9ld+u5ZO4e0Faomfk0G9mrWNZNq45t0Ew2oT+mzElQZXoSAShiNvjyxIX5KztjeWnpU4KeqmnaaU
7r+jaAmZCp/3PqO7tZ+F+/XlVcaLRizVnBwbYZczpGUnihrbG4BFwhugOqzJYx+L/fh7JPfwYum0
lbt9xQcqasq9EyUIevFJJ4l57RQhB1hRLHy2BxlcjDywACEPLXeBdn1UO7wYameIzXcpnc3jMi1y
qj2lircwbQiIQuUcRWLYjJaxYriz2syy1OK9pcy7rNB7zMn5eCip/GfdBcAS1zxsMgUsPOKdRe79
Bbdmh0hdf3/RSrdkO51CngV5BonydlFxIEuK/+BMorBBr1PXUR0bqch/NKPTlsAwrXgACyaO9UaW
GCGdDCg0sN9kVYmLzSWFZGIt3i4XNaezbL/KhGstUgbJgnaJziXOXH0DtZUywdwQuiboKdIX9iH0
LViV5s26E29WfLL/idSc9De8p+KZzjQEG/b85ZLEERAUF/93ejPLyDAaGOmHruxnNzWc3COUQWxh
pnHilsarymIwFxMbPbxXvq4jYvvaT4TdV/iOuMk08OeV+rrx8yKMlbsVfxw2wS+MPx0Bxfqk/xFr
WYC2OZLEcGMIgyABGodRCWyDuonjSdVrZDbiqvwx3FSgcIUNu6a3WdY+QumI1F60VBnRD/KRJ9NV
ymjG0RT5/9aT6l15A56ZSgMLIKyCC55J5XzR8BL3MDwkZdjc8QUKKbTmd0t0HA8Ru1l4nyqy+dP1
WZoQpFWf/PF/cVgT9Vu31SW/9CHdgGJbo8lt4AJU0dZyjfeEPkBaYg39TbgnVybWMItqfra7TMCp
yvnhYhvT7RoSkMFsU3tAWSv8qjx/e3wPifCsGD6kq0cwuOCnKSWYy9NiWiabgTwHW7iUptk0UyUk
ZOlRL5F7zbCkookOUW9ghnFchO/7EfSYKFdAlvhGiAg5lHqwi4FlUhsby30I29E+L3klla3VM7oZ
h3+11bKmZBMrm4eHPV5bj/BNi4504nPlH0xnid3Cq8ivq5iP8e6DjAVpvJ7NMukqttjmp2zAh1au
5sLYkOI5OPk3o9TJKViTTux2H1wTXh5HiwjlcQ1HQcNaC4D8JJT4SOPnxBSHp3IjpkvG3V8Hj9mU
fZvA45VlQ3Po7pjKydgcPDwzkfuGerkGvfHbVzGG9ivg1uQC3IG6zaVwtrH0xY3emRiV1rdRxQgl
oHoli6mkrnVrJ0kO624rVa4kw+1TJ36GNqnyoyDYbPxxcbDdMpRNk2+W+jMXGA/ljmbpW994c7qd
wQ/lpR9X8vbUh3p0S1K8hjHh7tq4CfBMgInjXH48Y8+DO/ioj3C4mbxn3phWS5Ro28qtxtOpP8Dj
vI0daKLW/G3tsGZkSscEhzDPOupeANTF+VDl41V3Js5GqCDLOrzQoMvJi9TdH/LZwEkDMIeL7W3M
Qqno90r2C69c4T7wLqeufoOFNsftAdoVa/JbHZB6AmVRfaNJCl1Y1BEjNQFkh2vdPPL42rdoOfx2
LKeBQjqkgAKoggluHTegXLg/qDUNY9c8J4PVteaUbaWtuVOqDXejJoGHWDh5egViu6+048Cp61rm
rlrWO35VUknLkNpl0sNZYhCkID+DJgzV25anyZy25tDY4p+9bCG7EfppIDfHrtdBVseM36poyg9x
D/Xrn9d92E74AQR1QDCPSFhk2FFT5mcYVsoAxVmOhmDlCAmVbqT/8vptSDIELd92pkBN5fcV5d4S
ak6W5gW6MOtDIhv6UEGNyBBlZHDoN9P/F3NP5oIZUMkXG3HjCgAMttsV4jsPDsldsMl9pArNovjJ
yhrBapqjQVi1tMSR0j6+7fnru4f3oRq0neNiIfE/uUwTTNB9KJVciOKvqTvlDtuvSbAJw4wKt4ZW
BKyYACBr0BztyiVEatFOvaF/bhmHWvgLQkdqfTkaWY0V9WtvlVsVGKs/Mekleb2Xiyf3+GxPsVWB
ZkecqZV4zZzBtmrssfvSbFa0/FWu5NsuBV/7dxhx5SiK+C2yrffwv52854nTn9rpY6v7aypGvpYh
U7bhtZ5G1D229vXGANjthD7G6cyWD0v6dmi5QlnNHzT5breqwbXJ3Tvi4C4G9/PoXYUmgxlVkSQY
99fWSyYnHF/y/0SjiMlk8H5FP6M6h/Y7bh/kdDxJzBQmLLPBeGkHmu5T1RS3lcjtb2b8Yiox9/Q7
Lyyk/OQwp2jYp4fGakTKnKzAvE80p+9WC2WWYsfg5PlBXjs2E1Vqmhhj2Vba/ZSUuo3XSAr5MEG0
lQ4MNvNpkpCWEkmoQNVWNlEYXNxHVeWrYc6U9+bIPHVGPxU+LEFXDSe6GeHzLMNtl1apqvCbKNE7
Jscs8xSvQP725c3+V7fAI6FrxHIUcA6+lPkv9DhhnOMAfSq9VaT0R/RShzHZJETwdAQmRPkPx8eX
cmBFkREbdxh3HiLVuwmzoTso5YwWV8Z4wpfA+TeilF/F/ZEORCEbWRKU8XSR/fwdXOMi58B5db/v
KBxuFdPH/rYwrm+EjPannDggYzhlinWEwyhlG6/ndecGZe/vlyusfge6daaTftDfgJmDdChFCvKr
lnn3B7sfk07SCEP8kKZQE4nagSBarYAMNRL362Mjs0oHYZBjPeJhv71foOarenNnB6XDbDtdRMxZ
daK6I+L7nzCNaMMpCxuNCTVhiZLxlDaFU8f9Rg/nuerZ7wayXEYrhbaiu0nKul6x54Cn0rRz3Su0
BKV3PK6GLAFPFUkiXtrqnUYBFnK/ODpzKYSGeBqqC6ansCV7vdEVIYBu2d7LCl9p9pIvJ1l47aQT
jJsUDAqNUsI5K27oIkdylXGpZATd2axFYBt+1++LNXtxV9GROvxjvBiSP3uoil0zCPe4DvCmAQYC
Sy7ZIpmAL3oyh9djJ9jsy6ra7Z7nlxajqjfRsH6rCc7Fn01eQbtW+RHyH9dxr7PUWD0JRvxN/Bjg
MPERCEDe6tjUwOfahnnXmnwJBica1IwwShKwI4eFTKICi5KmX1GstOk6HsV2jbhYOU98ezxtKhGj
XPLYDoa1QDtUXcIlgt6esCP8bMUqyUrzfdK3+Uc78PkbKjbnn7NBPheV19FTjVdwwQ6rH21N9sTr
nDdTNgc/5ARghQyd44fn/cpcsyGRS71AUzihZ/8t1BatN8fxfgAsxO/aoj0eyA3aylrPWA99q4WR
TXJzLdVk4YmQ2Nhml2N2URJ+xFnnYf1O61p9zcL1DkdCUGjCq59gC0B/+1s8mlW5Yq5FQkTmkTYi
nMrZjVq72a0myTz01jKCYemnI/EfugHBYMoggAWQ7CHxikW5kCmnvtzrSZLQqHPhokAGWQFLKbfL
QtFKRm6EhAH7NIQLDjFfOKyLmozNckFKWs5KEGZzyT0/e9w8/KZHCexGfu6qN2R0O/ET+qsx6/bj
QzPbBuihXXQKSevDo0BOhXA2lZQBh91uIe4rzLFs7Sk5XkkFGeSEYuiJL+N5QVAMA+RB8aSBLYBk
NhYAd64q10HmIKr9yhSRg6661o54cuHuhW8xfOsNDouueA/f1VuNjglaMCZptiWVIhNVJXylyMth
OtVhRH+Tr5+SDe/Q26RtHAbjrWj1QhXOs6y9FTzTl3vEQDbyXfuHPnNFi5REbqxj7rlZSUm6M4tK
XKqMFz+v+X2QidyhotZ5wMbeopslEIlQd3HvrigTj3LA6HSGOLvTljQEPOa9XYi2aUftkVbjsWcJ
g0LGdFbPrmiWgJAIweQFq+K+50ckqqZhrO6wNP9FiBnLpJlfn/4f4l6zyU4uv03CAOR+HgpSQu7P
0AO3zJQB0IlFZgycqEFU35LM7wH5kizZBwqhTep1LpNBsqqMtyFmOqbQneT0SGhOUUNYJ13K70Tm
BxfE24VnxG+SjivM/m9an15UPE+ps86T71bfKEan/DxQNQvYS2d0KPD6C6Umm1ywmwIyAjDOmxY2
XcAOFcMsNq9g+2uCdihjU85FvNiSk4qRJagO4wAg5ynaQuiCladGTz91g+kRu6YQa/RGuJhBZBRu
KqLeFQLG8E4nvr/bfS+UxBEXAfiOrikUEgl/zhvutXVB9G2v1oo39RZlHSq04K16VGmVAi7twfjd
EiQBl8mk37rQbKKTHpI+C1pjzQPlWjJqgVovq9/otIs2oVnncjgo9IT8XvLvBcKIry76AdnyFf02
g/c9hiVvGjUJQiXbY2JmWhMqrpFTEzEw57JODQ0puZGadynsjDarLTp69sQKuKh7HvRcJQ/psFZ+
QGHimgLOEOp51Ngy77HOiXS+sBW/ydGyGfkqi1NsP9SMdY0999Wufg2hAUvY2ecY8QOXvdGD07wZ
ZRkneKf16+vxxjUCavG64pv+KNkri0rW1SIxDyoZmtDGjsVXe9nMlehcvpLpcTuhIwiQs7ag4Ips
7zjZyRzXDDzTi9DaEpsKjwhf/6AsKC+XUbjzwYjI2W1gBLiLFoTzgj/ypFccsBC2cAwT4BWptvhE
WvEQWNzoE+4CTPVIKlCrIhy7THlJe5E+Bu8JBhA1xojkEo/N+1SsoJJ+3gqNJWi7UuqptVNv3mqj
yVtI6tizKZMRQgMEiyofluls/ERMLVQHKWvuKT6Q/Z+sEU68nLRH/8Q1DiMnRnWA2tS4oZ+5bg3x
pJTRkEm5Ij/KP0Ld8oVoFpljjAdWoBSPaD42k4KggKZB0Py2W8vRlkFVwtxYPFNZqUvMn8c6zWq4
DDFo9k93BGXPz/hHROR+jrjlAJ6VDx/Pdgv5LSpTFJIIUnTB5gSL+SbWFj1TjPD4Z1kuBLtnWzWS
Swmz1r0vI6jLdIMeV8cFrv/v53bEWtsLhvSnXvsEYzibsaLz2PueeSfc0P6vQMhFOIndXo5VER4d
cs8cPrICq0Y5yZugLOH3nUO0WuTYiYQKulSUFAMj1GDogMT1nLCeH2f0sOTDEPzTntJcfiRJOKxs
2DYOGNtZYcne5wTso7jv5pJkHDnuxXkDSk7YhywM9IbD4tusgF27eoLzUIbrpXfZ2j2g27gClh0c
26cXUURgVlXHuy8czXImYm1eMB3tjuz4A6TUBUmm9Se8wB8JkB53KY+yJRhwW/9JM+hYW34z+Qti
AQOOhFOWRm2z1a5DC2uf7M0h6O2HNF+8oj6BuGSZF3gekyoXLTfYYff/ghYMG55q6fTIPo8jS9uR
ixx9PNRvUIbhgaoCOqEmhy32oUp6z0YlLMUuFTkJGacOiFh0Qbnw9lZ9f8AlCETK62o3Lt6hHfGo
hOcO/khDoE530q4GEuc0RqHkLUZUhRgV6ulSZZusxeLr3/LdIST0Tl10RQayuzXa6xpTxH6JWCtD
xEUd10sIq8B+gkK1i7uEOX3L4tbCv4WJ3pBV/B3HDjHniGCRgM90rNlnPlbgBywvGvHTdIlCEPYV
MqjT47Fj+563DA1xnr7D8P5jHXoySKtxb43mAva0IOMZC7NGMx86lh56ZfsCnQNXmzeGS5Z5E+Ak
df8i97WrSQcYFCdZd9SUL2GpMg9JykA0W/4j78kc2deiwcAcIizTP1HYTgUkCZ8QIazjdFOrcnkz
2R10hPLThY2nLET9gxwX4PK3QGSO5yFU8xYFZLzrObftcNmTsy4rWxEoxXgMQK/duyXaK760dhJX
WiriF5QegIYU2bdvW9jh+JmxVNn9A72znoiuV/l+WJR58H6nWZSKgxcckJJnbGrGdX7xE31n29N6
vLCTE2OU3hogQOhiSFk77dROB/YED5zUyy+xUohnFhcck3U3bRtp4gIzr5Kvv9AngdMoOt485Gxa
YBzs78T0RcmJoWPmvhVPGuxoGyhfUdyiZLnei0x9hgYTz6TTvZSyTLrGzxyyDone6uN8e05PVNgj
Cx5PN7jAc39zOssQwzR7HIOOoQf01mIScrE2e8t6Jq1+OzcTYQARnaoSBPHzM4U37gUJyWMk/cvl
xIFgmA8XuO4yPum1GXyFUVJ+J3LFAfSAtGof5CeHYAEGQenOY0Nyel06xIuFxbJmuAGE8rDFphqK
VJFAQeeag1Q3mn13UVVjCv1D9oZ0CYTb9D2SlBuNueFCcHtm7VpQnuVFk4zkY9V49cfwEXhVEMpe
e5O2cyR9CR5nzuwZsjXNcH1NijmBEzuQpF31tVzzXekM2Kq7P4idQZOd4dlKFKvEw9AnSS4My64C
7UiCCPoLK43eWbeWo+smfvHuX4xxx1tp7hs5qUVlvVpEwzBxTzT2LSTJqo0JrXNAKYvTP5LKlsRM
/Ir77WENtmU6VncDBLQQzuSU/daZ4SXFG3Vkp1RvsMOEgxEWzmyvbEnzAbrYP6Up5U9R/XJo7ym3
k0C0QFkoLOerpp5pIlUi8rtLbmWvR42xDK9+AwSe8xuihFP0VxYSJRlBhioh0vEs4H2wGS1lf2lE
tlzvGqIo5Jxgr6mrrVPbBHN6T+7Ktkf5HT02dGgRvX90INAZb+KScPLuc3zRW8X3BkApDKp2x/Sc
X6YcDzKRYHU2acn/9zOACQiLNElE1veps4/qlnLPd9ddmyXstaLrBeVJDgmkcrWcSgh6vq/nVXfS
8WiCct4160MV+B355JhNmTudMJhIMU2inuVtzcrR1T3wj0jziBzaTTf27gFLp2/ADRowBdSWoXiA
EkTlwVxkv/Xm1PCnsUgmvIorAjSQnywKYF0psm6wkNSzQWP3Y0Dp2F5zpG51idRLaHss8md5m+A1
Bzu2acLQKvgdw0rWkhJ1w6j3n4AtpcJbCcJvWdwXxVqoePoJ4QUHdGD3+przmLjj6HhcH8EaxP4s
kZicP7qmb3ROg+uYQrujbqwNUUqiu5zBBc8uFemeYZ/4ChazdMyUs5Zmtx4KPQxOTPSaidRHGTe/
88PdEqgdNUcZPQKOOEweKsN9VhEwKfTnJjgIplEMzM1HHy/BxNZIAPzl1HIjyTfUUI0DJxbNAN7p
0VeecExThzGgtrdf1WVyuYbvxfngC9+JvzD2Q22ArGf/Kt5yCv9sY/6/JRpDWxNp65hPHzfR4Hba
/FUiwlt+B2gJa2k3mV0gKLaZDh6aF66gmRnEf4f7BEMtLe8S5c0WxQ0e9TiidSFVtm9wDSYsxH0B
4pEVXYSIKc62cpeyo6EIUcwxZszFZQMsRGkycl9yzMj9uLFoTGzjUuNcg28/SQTw71xBbOAJmEFE
tqtvu2YUHO6aOlOwUv1+Z5QeMaMKN4cIMiBccfKHImjTXYJRayf3eLSf6zKwE8iYa+IC8e81qdAc
AHWnWqQ72cyPQPgOptxlcvvrGxzWevUqCcBww2LGd9dYAOYyXHdqS/4rYqh/bM1ntw2xqKi+v4DF
SEVTMmC/jh33CKT1GwswipH2+XrPRgIENo56msBE/iTz+lrujVJsTTCtCrk2tDzZNlBgs9idi4tb
kvSOR3u/WhUtXheXKJ8n+bKlWsmQjWsdoPNn56BH3xlrDUtpxMD6UQcZYyT6xZId5vqxF+EPqDCC
9VvzKcyivP5CVQwBKdav6DrMqc82EniRKTSnCUIRzhiI9CYWq9HbwWZ/q5lbS2iUMqJmGgbIuGjO
cRiZLzCxBWB6zhguwYDUBeOlZt2Vhq2sKgq1I4Rk08BPjcidzhrsmcBVKy2oCLEnGpKlvxKGVnqK
6dnzcWhossdhcP1XrSjZpsLZwgfjdkT9KxgMH58DbIi7eg5QWTcsfWLAH9pPEIwwifIuiKx4WJNp
9i/KHIRHjG+u6yBw60A+MlzMqv4r3O0WhRfiFuDhxA4XOJReOJLIKC2MpE2hEUO7kbdMRwhWVW21
Bw7UOW80akHTLXAJp46qPIpybGyLnvZrRrE/EMp97m9wTNWrs9E7rW8WMD2ByTOwyOl+blXuwuZW
RgsADpOSGWFzUuXwmgRQ3qcO3LzY4ky4+jOFSbZro7I5waClYZO1IMMr2aCP7khJKGr/KhRiBSzT
RaSvjAAnj1afUWdhVxMPgtjqW7ogwtWI5GxA4BJhcR1XmJCys/9EONFc/mXbxdoltLQPKgusUvCY
75g41wXpwELRpziwCGCJTF801HULEn2rMs9pNJZPbdbRgUc7GlXMbd3mX3onLyzRxswdNMz64+UP
T9WxNwmXHoDjDFyOyLu9BWILPOQ60N9SGvxrET0bm3a0p+eGG2B6I1T+LpBxk3s3S5spVccdQcxs
K38dKmE8tgpf7qX4VYJ8bEiT6AUye2QWq+AKzMEPHAr6ZdysTW0JshOf+LNEREyUSjvpXO/cX7fj
xfnZ7UopeIsi6jiYBqVt1/Wk8fnDawK6zZUB6cHMBgeoF4zMxO2nWdXCoUtVPCsBrkP5Srfl8hGS
PMVunfHkUuAxdv4Uj/DWt7pQGBjQNKpgTZvpZqZNf0kSC+hXlbPQpJMcY60gvsUEKkNZLYVnW08S
RQGyS66ZWroW46uX+Q+LQnDEWgMM/4ABfJamHUncUomUFBg4HwLBogRqHTM/JE96PF96SpqKXepU
kJQS3hQhcB29JdtNK/Z/0OdqrAlodX4XpaFHIlsWO9m2Gkki1saeLJjRkAAa+lmtIzCPAZnkEIwQ
jVDmJc8gGda7JD2/KKw2xhHpG4GltqnBTqFM7QCS1u2xir+IbbKSeoXjg2okCVFv1rQVILKmOofE
DZwC6prLNFtIsc5tooTqlFMUiDBXirnjsyrEXSttRsp91rTxSARU69FxXbLkJ4ljGEJyDE53djHS
+vZejV+unT3hHZCXhrTb7y6rfL2cSnxS0dP1N9cSIPpES9XKINKsFxBtrMfo+AmdRKGxZ8lfLkeH
oRYdJTXGWt84mTrNKa7NdJ1z4Oyylq1Hk1tDa4XOv05vQTuyK+rFeUmJ2PbtDUBUquf3OxFeSkwN
1HjGOP4vqkDUi/OYdrlZcp99M7mu2vMhlyubDNsTpcPdYa4pzrT0NTpNz0yBrBGQDPbBSmdp/XCX
aDWF+tUlk5TO3KyKQ8qX5B/sdL+CMie7VbN2KRR80RdI113gxMTfuKPGwc1HaoLHybeRqD0SgkDC
WD+eLujL7T7fDJdfHqqQr9wJUTxqBcT8V6479TksZrw+TZxO37Deus6pQ2YamhgksY6IEhOLZ3sE
8EhKdVar69cMYg28/5hLLJsAUJVZTD9dGyUDbKJtWrmQCLQtWDbTDcACX3m3QqnEWJoetwt6Sjv+
0tCE6M3AJo/jDA6BaPMVpjlvvdklribImh/C6G+Qw50fYfdba3GPQmDVdzWAjvTK0k1JQAPE7+rC
Rk0eqm+JLqwcAs149aRzim/x/tQd/d7K1mIKzcWemDq1Gymvu0SQ5pdvJL6xylFrMSRq7QJTwLeT
rw3sdvK+04aGCSsAEstKDWXRPFQoTnD9k6EZ8iMCpNmar9VcoAkPESFtsImjyP1qKuTooeRasjlH
DSGl1dMDrYrtsA4FBgmdrQCsgXikhFBHXQaiQJj2xeOxEG1k1EgXebpiIrqSGMHGPSccvwTMX6WI
l9WQt4ucnUeYa1C4D95s0azirJeqjbjCSK2Fyfx7S8pzvURz/DS2VVc90+umyTi7qosbzFB7aUJP
qV8wMononjVEs9AQAxzHORutBBcTEnwPnonsb6kX8afjJynHKHzXruHNFzI5T15A2IwuES3toE9Z
vERxG9bKcRjZgy/QDWK4hPhK4OciEUNYwzCWKXYskkT92/rN1UCZmxApbo+Vgn5iMeo39Th5yPaT
plxHDRgpnF1X8s21V6fQuNH4gUU+RS1vLQh7xr/qZmVmSPlPwGS50Gzd9abeIjuMiw8E9lfgAWEp
RrWIDJezznXw1Y+JXZhOdfMdbUVFr4uRurFBtC92qJKX+mRs+aFbZB5DxlHtMdN2EZ6JGF3RwIkD
6OqU41Rr2WyArrtN26QKV05FHJdA4c7t8Vg9De5iq2oo0wG7Dbeh4eGSsK+zg82pnJT6hakTOqs6
tra+5Fc11TN0T8FxJIG9jSekVRkZ11tFoxs19KL41yni5NHpEUPoMy7vgFpvgHN7I8L4ThC8V4Tx
ZdYbpvzYfM4Y8UwC11PWgDoBQuNQfvu8Bj+fNo6c1mGavJdXSEDUErS1yKTFiynE4p448uN/Hqjx
aj3AOHM2qSETfpdVJ9nUcFWimCVzADwiSKys2QrvS9RYiFbiVvQ3ytXvsrGIeAoK36uu8GyimUM6
OwfCIK6MiWH54Iauv6eEcv4WI0ulC7BmQjXfeB6dpDMRFESp2salYp9Xv9urBIKzp45nf3Fz8AQ1
VgXRcYygMJgWwiCfFYLkhpdmSI2BPitN39GkUPM6kYo+bpSRekTipjiFcba/o6OuTgnGrqQW77r0
w5OJxu6tf/5tChWpZEr6fbPyk7qDHkGUUkmzfoKbBGOGqqQ/UXuhzXVzAZmuKlIqu/qNcUmQlGTm
E2jE88kJC6bzHWi+q52e98WolzHBlNRcEguuuzU0l6RSGjYI41hv4Oboquknkvz//f0Ln+8LbOiz
XkCkOTWPUOXlWWH38j1XRksrnV9DIfnTtKzzzMpPU0Pm5+Wreme8eFGL0SV+kf/+bNDfYWLZnSbq
zm150CO1MKWEY2VuBbnu+1kTleKY8cddiBjkh4VrznqZzMKebadj73Se9keRKdw6U0hEklZ0KLfb
ogn7t28wyS2UwXlDwkbeWa0DbBCBPAgcYPXslLY5nHEBdufLT4uDMFy3nR0jJKH2Y0kLPZHUJOBc
sD70ELFEdQ7bp3Py6/xddozmIOnqoxoX4dvfRwF5vPBIX7M7+I+zPsGlW971HengETlmUyUIXD+V
o+DlmzZMmofFCrJpuRJj1y9TE3+wPg1/ZymJ7drrWvM29YWqfC5U5ze1lhwDi5WU+d5+ILmRXFzN
MvUR084it4BxnxtIoCU7qsKRRMprhTNHKHWGqj+YGgwjRMvuCipihG6OmVWHnT3WENi7hS9R79DO
Y0qiTaK4MoRYLbZ3o1b9aNI8lZIVywhiVYHgWLvIWU2pv250fXjELX/cB54fmZFnvEpaH+IZF4aE
Ive3CcDq0ufUlg6jqkycYVpQBaV6n4InKfiU3NLXNACXWhv/dnQBCraE+ONJ/pmqLb9GHtH3vddp
XwSS4Zsni71dE67E9embcqKx+8foTHHGMFtveP6x5oC9NYfr0y/WHR8j51bOkyC5Lv2oZ27eKCPY
7zaVOdjcTEo+77zgOYPyqVi3DYVt8QvZ+dfOM7oyxvfawB823YAzYCWh8Txo9A68xEJfgfbK31g/
FXjYj2FBPqVHPF3WqOW1yYTI8FLvEWnnZwTIyOa9Rml+XMbEJ0cgAZkVAb5tKAF4o7DZTBJGj4Hu
4gr7xMypnwhX1NLPDOqQH5+veF/Y4sjBoJG2zN+ts/rK6cXB5xPQZ99zEJXtfOjymoKi48WJBnLk
nW8Cn5X7TnE2i1A57hmCOMNEOkJHgD6EZkA78q5z24AGFk/OivOrJI2Jt2RhExun9xaZvILvXtl1
sbCZpb0tjK0YcOwmCVkiNsFk7/Nhc3n1XEi25ZLcPuA970xZpYCcefMcnr6p2VVh6lfJ/xdMFocZ
8p9LM6zIAm75Ov2NR51/PotazZBFzOAgLVqMA5WF2+8KuEp879F63JRMuth9AltR3O2Abiqxq/b9
P+Af0/ZYahQSKgRbnDANN/xHKcgikeA3kfRIkfL/WrK3co4cu8ELCgSg8UTmogriaJuUckD699nl
RTFbW7zuCbqIPYm37UzRWD77CPmlgbv+109Rw7/l5XV4qKYkWKpAYoJfb0PwH0nU1Pib4AyRIxH9
No2H9H2SzB8kDCa5ra0C3GEmr0d0+wjOBflWcwGdxMUPXuq1ETOKseuK9QH5PflvD33whElzsC7o
/8psmobp8J0eW4MMWxZM40tsZrm1hRpRXSb9cdop9SUYNCbuIZrsQOSr6PEN+bUTx2WTp9yVTPES
1uJRgfqmMNL/CySIxnVQPgSp6En2qYxzNdygqb8Nk14h3f52zAkkCZtUdrRdFg0ved6Yy3PSYlE4
3NPfCF15y2PLDDSOEXowL4P0s5xGJUEk3CT/LF1LzxdqADXsd99gUM07z1cNtyqhwPK9y4MQnvwf
HqfyWcXFHcj/Lz4z2nMb+jzOQbZR8oGTyd3ChAwqJedTiY6G/qT6QUefRjrA1cFF89bxYHHPAqWg
Qpof2cDPcOBwdbh2gEwa8NzAGGoovCl3ITv5bHtUnIOoAcJusSxGMlU+OJNAIiNzjf2SNG7cWOF3
2YUJLZ8MbbXXNsiODG83QtSSJAtCGQMPQaDFBnztmQmDv9af9oP3LAuYgUN1Rxr09QoBwXywOlES
g/Levza0jCYF6XBE8Lz4Y25v3ScaMmHkD+YkDnvFQgYNA/iRqN4+nddWKjqS5xKC3RRho8gDSvy5
FlT4k/DH2lnX3b4hImdldxVPGsEnJ8LBNMO/oKdJCWuixTRkK1v9hF/GkU5Gxdw5VKnHW7AdjWMn
LWaqchVLwb6h51OZyRfCIA9X6ASLX7AawbYgSy8pGMmOggLHZc6SS6ncTx/37oeNljOYgej2S7z1
JDpUKf4fj6b6348rBROtOS7OUsOU7MXZPr5vkjU9P1OSZgij2GZaWnVa2koHnOZTLhAtmKPmuZ1k
vrPEBZV8Jc69dmAcN3T06Cp0hztFF6acsS4E+bpWBLBRkXwM6IA7mkgXVOjf1xlYwqEzI3tLdpmF
vrNsOsS1Wk4ZvAkA7Nv7NSFlsUyV8BdUvwYEaPParTZxRDMNkGf2kfmM+QRrcH7ZehhgiHApehQK
/5PMaTf3QktkhiiZ6bQddh+64GxxtoGffxa5J/bdBC7yYG32F4KI7SLM3uQ4XLCmPd64WfHcYtMq
ZsZq9gL65jNZ86ZcCKdMwdfoYaWevFjf06My0w3jijUA13BJMz5KpPotdu61VbTvLOs7K5Cy5uVj
2xekWCjJfJYwMFAS+tj+xQo+TqX70PkJFcmF/q9kKsOM7xN7IxyIH5tpLxqLMR/NN5OeJsBGjXuc
3q7l2fvkZ5R01evPbEfApASVC5ARtJEFif4KJ5OYt+I+UONJgtJbXoZ91H70aGU/dAeOjj/r7qCR
Lo3RAGEJtQlJVpaPexBpwjDgWMHIEMYlsOQWTD2TSQ0b3MlVcu/hm205VUeaPfQBzupkTh2p/G2R
CdY8n9X4OSuUFS7Xflqlj8bvGBGbZIVibz3K+uCa1/npXLkAIikop6S938/jgOzzeHSN2c08VEfh
gStfc7ibZgoC/SfKjllRtJk+/oUyHmKlRaH+GNoqW1akKRbw15Tfj6nb+n/h3zmKEporYXixipSS
xgxleyX3M9CcZjRhKGuZLdcplwswLiBh0MX4s8iu5dlIyXlVNYVUM8R4x00ifAO1nXDqcSbmlGSP
SxsLoi86PA4FxHvezuYZW4xtQp/on5UrILCavINTWw4dhzc+EsnoItOTiPWyOH5Uypr7DgI/r6NP
VGrlTO426umCNXZSc93s2A61SUfG6q+nrpMsmJgwTDsbNxUDLNXc0M/PtE9dzgA0QvtTzvKkduOL
Irp2wLR+W/jAlm8PNU3QbzKwC7vDUuTJFUwn1AFQ97ZnyIbyE69BA8lKWj8CPgSlXkyN6SXsM+y4
JsJ8/IS/JRFWhq58ps4OItkZutF3yELqgUmod69u1K8qIHoyxbAg9RoqkPCtH1tZ7gppaEV2H7Ed
OVfv3cb43uyMnUa0hqphPINk0/xlIyU02E7N00OUL1ogGcZLJQxZpe9fV/rC5U/fGrHlGUj1K0zR
5Oyhj1ayPsfIaOCa7uTOItqgUNM7HDrAEig3QAguXmOe6PG3S+0q2hTeU2Ikq8P98c5ICNOpa6sb
IHnmdWrrITYL8g8+7AjegVxxuyW5oZrX7oW2yEXQzZzEbd6oMeeumk0Qbf3zmeuaioA7doljxMx2
NwZy5VBoV8+GZCKStkCMKeTzUxPGr9ryxxWHdyTsHUa0+DtYFD2UDmDfaT0PYZHGqz5CBnuQxpW9
/tLj8vaCAEVoc+Y9HAqxWrFb6aktfXb3HElstvPnvUK8tvOfslRhsYH7n3vPQd4vzvq2zBl11KDh
tUoo/ojv2AQLMAVv9Kh5ow+Q8bs78EqsmMDV8+SOw1MeH7qO+6pX9WvvU62M97gHiTtw5r8+n8et
kT2BqQTHMO82eMQeIxVKfmMKTfSUedyJxEe1ySvB02K9ZeZvJwSquoHMpNBn2fpYBp0fKRR7hqPY
SRFENNQDIu7z6pCc8oIR406TLJVXGV0JGhd10tApmMjWACW2sB4MH8b1/l4gVj8oMlFqZG3niXwt
FWJGJE0tRwMoQeZoNQ0QqVUFKRvFQy9Pu/4E+JKK1RHacKl0CjgZy5TqVIaw9rGGWkmB+8MvabK7
VWuagDdB2rfNs1WJTiseFAo48Bnh4IbweBZNsXbbEfG+o6MOXqFrEGAQutIkyBR3owIF3VqS2Niu
RSKfdiXep1FTwTfTt8bvMI8VaKspI8QZU6jaOPOUIShOZXXfPpWEcueeMdU0WvJgRH3cDp1C5Dz2
pAHimOtXc10vt6x3gYBSdsGB19WrkCSxY/76VJLt4uepG1hsIpKsG0Rm+ZOvK8Mh1rfgrPI7aA5E
lkA+/KiDDlGI+zfLhK5KaBnfJ9MEyzTtIl61q2MG9/PkEj8oSJ77JOMrHIC9Yjg0GSkpkq1Coh05
Lcd19rMLZ576UGDLy8/60eofHJrorbRi1Ur+ZgL82+75Y/D7ccPuCzHx++hSBDQnsTWgwHiRnAst
3GgtXiAowhpHGthbfzQf5uYadl4kbEvC8IkQ4lI0JFghKh4Y7DODy/CCHMJOsMWDDiq2FUYndUAL
BoD0taQi17bfGp6Eyc64l83ebQueyjCcDtJHahrmMzjanPY213pGQAx3sqjpJbMwJHPPi3qFsgu7
plQpw9p5gUyl4cWEjaoTlYc6Vg9XIVh8OvJ6G4a3CAGZz2vE4G0k+axJEJNoqU6Q+/mZrwvtRkru
7Dl9UvWOETa2OpCvtWMln8/VVKLlxkHhEJmAgHwK9z3Ck5MMEcxeGJKwpvjVuUPzjcUPTOUCAPC6
Re05bBybC+Tvc+ry76kjQw4hnlgbz2F3i92jIAudVlcV6sO9Px/WRmf8xVXuEyYbnp3MYEt2B0lu
TUV/9UqPQFAU/yG2i0yB/CpOPehmKfBgyCm9/TfCNxK10/72OY5fxPUm1vKuNXlAbr9q7nL676RN
aXQCHCKtg2ftW21h0Bngi9lQy+tqxPRFe4o6cmHgBHyNbDoW/aQ5NpcsgUcVe3sFbYNvF+3Em+Mh
r9ujUMqss0y8T/H+5gFPVw5iUxy89EFY98F8BHYbMEPSzK6Ht1cd227G7npEG4RFLbs/xUHgcWLJ
15dQjCG9G7L3cAZkdlyAiiNIdiudp+4pZB4yp2wBZpzhuvwS8Y1slbfk2P4qtUK1f8+8o3ky7P97
FDZXXcD8yEeaUjonkvr9Wv8o2qMHqKSno1YBsG39DA2Z/q9/GzQyYPHO+5LwSAtyymY6WtiP/xEU
bvoJ8REQDPX61ZShqq4yC4YisRqz0gkZRSZUrnN7jiUkjPb3GOQZyXdKg4NVVDd7zwR7CmyyKQlT
6Sz5CHwJMwK8EcS+euAdo60gSLJYb88CzLuhx+avpsPIzpO00PxpSOH5T3pKV/opnuHwbjL6w6Ti
ykUl3ul28FAibJbU4dokpTWU3fbNAX4vL18r1JgS2KoATXe/2AQhxpC5ZakqO6zsYgtDcdVCy5XV
PqwrJwOLO35tGYfK+AMCan5Y+UnimqWzKmdQ9O33oyKSCdbIVTzhkFxHUyHJ+6K4RV+F86cz7mte
2ou2sDuPi7cB+AokTTkgjMhISm0s7xv2Tk80Jk0GZplL4djRIQRz3PQgDCFIn2+0nxGLCRKp653z
zQlEK413mcvOl637H+vIbBkgLtxFhoiitMwrCRmk3yhSnF8U4psqpQcc1XwAkMCHh9PuI6Sr651o
DSVQw41ltlif+tbnp5bjFfERDgqnBMpHVcbizIz/ZNfQmiIueqzRqvPL2AOHOTKxmdIzYl2hzC6B
r65BA6KcL7/zcr2UE6RhGCYseDcf380VZyIb6mPrYVADsk+M3FkMGEdu5V6amN5zbE5Vgt1/8zSN
dZ5g9g53YlmW059WhQXEimD0wbcPVClt8bF78O1Cku0fLEqATrIHklu4aRk6X7XxGmNiHoKWNg58
6pZwkpCvdKShorxeJpI52+p3vgfUFWpqbO8SqhUXkNfDP96SofMdkEfEDgubmABRSohtewTDpTiQ
qpsJo6sgNkYyk/3N1GmySFziVZVDtwA3buGmKCNtY8RAxwbOpCVsc//YFfX5uLxWR1aFdFza8iuj
KkuBi/eLWktzqaRrcPa1+gX+66+OSsKHkvDgWXb66vklok1fcsRISL393HTb91FlaMf8uDEbiA9d
7eCBIvzuAZkM6/1TdZ9Nwi9wlzdvipxkE4p5zCLrtDSUAEiWLs70oqHWi4bdj9KFULpsonPIpDyZ
S5Zw1jMUUYexzP1DBy+tIkClmXNTGYAofOpQZARio5nIvGzHBVpJdlCTaVzlMnydpGrDLApvu5r6
Kh2+p/iXAvSYdiCzm2TTAadHGz6VIM7aN58X4LFcdSaT/M52jXyD98157S7okFO+MFKXdSDfMtAL
9sJQbX/SUOmJ14fJnOc39svlGXMjd64r2g+peoZvdcnl4L4CxhVY84eb0HftkOL8dj6Z5+p+vY2T
MQzlBZ0qr3ceQkmZWzso5NHojwyC2eBu6a5ZpEMQm43L9l6crJHT1kI0cDoLO9VD2q+9G1SdM/pb
FLRMQUhBV9cHQCUTz9DHsVXztswU2z8s5s0jt0V4wqJHI9rq+lDywrKF3nnHh7tSVjesgECgDAmq
G68iXtmoA+lEN8C3aAIr5mRWk4s5lbQxqiDXzAri5b0v5pKXZZzq5PCiKD0vzeQtbvn3sgbtJJlA
xBbGJCuKZsuSt163xodsbw7YduBT4o5snOpRutIQ4yylS7js3X7rWhiyEacI0Xpv4hqrQNAxzu9G
BXylsRwDzmf3JWXojt87qGPd2y4FN4EOSKnvq1QFW0xCgKqrfw9MU2EyKmcy770e3agfAGoYbUtu
Al3eAhsIrEhbPH901YsM/5P1ahPq7ap9zWua9vVZ7QIkWnydR0maQ57mlzAmS8A1VrJ3sM7n2w/8
HWXx2kkzmjOaCBEzbWRGp5CRJPx1gLNpvRIWztVUtsjln11nk0EmTEGu5ig+VR6K+yp/SP9XwMlg
ZrAOCKVZnLf2KkRWfVTA1HoP9lwgB4HYENwBVMutlyaUEstEw58YU5jUL3opw8YYgvhB/Jq8GYvA
pk7X2K9IrRarjZXojB1qYau+sGgBKgJfhWovgYRx4xya8PnxqEbJLOp6Yn+qeoyIlOfRHwpvAKOP
G0z2M6JkA/A6nIXqElZSPjJiLaWpLOcRSSScaz0SVGqb6NM7uA5U9V7aH84BXRTkJZX3xeXxJWa4
HyiBImLYd8io5fG5V/upNZYOsaqxONq0sYUzBbqih5hbrB5iAqj5PTQukPreE+6mXM3VlbJLHIm9
aKHXkjWY9eZTpJcPiTCd+c3K5+yo6wSngJo3xsE5YJ96HVhshIrmQNZG48j3j6Ob1a5fZS88ZPej
WIl+UhjENeDdJ/vLZwwHMiE8UdIkAriZVwiBeXQGMqnkPDt6lxaaZ4cjY/3RZWKcj3ECMu/rX/b5
FaNF1BrrC8ATc98FKBEg7UHworrnAqd+sKAijf6mjwx9RiBec5UnIWAbxFaj6THg48cSzBPl7Ta9
+BXNIuZ/1imC+dkffGsJgZxwhiZfFvJ9ew+sRjmnp6GWoMB8Gx6w7moNtOrUezSSelkstTnkjVGU
Ej2ogzviXylZtKRxBjF8EU7IOJrtaCzs4B3B8Ab+4szJY642s6pG65SpMFQimhottsnkMZaoS5B/
YHeEZ2cLIPWVKqPsQ+QFFlggXC/zj6r3eNFaPecl3C7gJ2mCzzuifWg6b9/R/gHpVX9+anS56nw2
6S3gyPVXyblfW74gC4DxnSowmp1t4PTksy0XIAJx7cCjN7L9hNnZEoWGO7yVJDu6iUjjbAkuFuVD
q+hBtQIVoyAyB4FU+4PoG7i8bVPtWafnGSQDpZVnPtzlNTJVhsB0YJm4z/x53NqxMP9KX/v7kULS
07+ouiaY5o4tf2hvohe9lChxi6D7IcU5/8K4DHogoOUi01pouFh2b7hkantAQtRpBRqAe68ls1zr
0WDYrTspotYxONE2qpQvubqcdKvd2k8yyCv8cfrfyRttXXOU3cAU12tqqJi1uIZAW5NOfYQiUAQr
+M7H2npuLRP40nw5kDXhpGmvbFGemXtGj7sU8ck4k/Z4DKp67KmolEAnJX0/X1DHwXhU5qPXhNCW
YceLhtLkgIiow3q8KTFJrzzYKMeogZhV84qoSJQYywnla35FZwn8DYrYjy6qQAS8QtJcNilL09VU
xaMw4sLldS1V9qmGMlZ4tsDPZhLcw7Rqt142nZG8HgQBcJkPFhsO/TL/npSKNkzaW0QHHWo9S8g5
AMTZkyzdrKOXey4EVDCS4oKpPhzo1VfIv8EM3GTADQnlZ1PwyrZWsTOvVUufTy9rg02t23M2J/5o
LJc9zvgoL86bDp9M8joWFJYHyr04HxzGhLnfGGSmwfjWkGOUdo8jQVq7wn7gPuXPr8mALzyU3CWa
J3DRVHmr9vAnMHkBwGmIfXB+MJXIiU5C8Pt9zd295CXy0cfZWp5vyIKKKtJbCpFGoMcqhsq740m/
m6vYeEIiBGp/5zhNEX+vHbCWfAkT/CXsAJ59L8bYv30P9RT+ZoQbeC7EFfSPNDznpbPRpw60ei8A
Duf9gY8VBPQ4U5om775RLtz3VK9mCh19QG9vqLDSDPbROVmX7np/ZlDfdIwS2OLInWWwzGMTY1oV
O0l0ClyTi/H++FLq4fvftjwDNgyBAZNIoU5NI3ybw5V0bW8uZe9xQrTcWMAtGsatlDxyRAyFpeEM
wh735XPJ6Hr/R63N0V49Vuo8Y2T4On82XvwtHysRR6Zi9odBhJha8qGSd/KrEgTQazSiUyqxpjgG
M8ITBSYoFpoiKmogwXUmYmhRX0IXCkhQMVda75nrltU9B5gffvOoiEZ7yAt2cEPilCZUUPAcs6GY
0nzqs3h+cgBQX9wbFYXyagIDtlw7IyaAuWuOCyMhbTS07+Qboxvwe2ztu6FJo4i9CAxyGFL+AoS+
2avu/Lv1V2cbUaIvON3Vdwv1enHG8VsURJEzF08kSmJA+J2di8N1jtZyQIK+KuHXyPK1e8Y8coDv
7eSIwSfx7XQqDv5CGYQ70VVsgGjRhA/hNzMr/yjv6SeslamKaIs5vY+TKQu9AZgofdfdPx+lRSm0
NhJtDQjCbMMpwwNKCai6DL06zEqoItLTSPW39UW5qyyN97BTutKxgDt3Y9bCQkpOw9iXmv2Johjx
bUabyvkIsdoJKO8ImHuef201UhjrQZMdT9/JY6uKfJUZv8/U+XwW+JYXlj8OQbLglwVKlIolt2bQ
Dbu0ire6kzdFRodAwFgtd+TmYqYtWghtukPZZDKL1h4OFrR7qMt+mIIJfT0z/1OgeaOv5UAODFuo
ooAEpdimG92O7H+c/hxZ/rtu48cBSyiLrCtMUkAqELTPnA9FVifFfQTgxmPARfK0rtrVtPLWo7tt
ryBvrg1n00hv1D3sqm0X3fXbRHAB+K80x2GXrXfFahh3WmNRZxl4akgrcgc4TcprB1Vwv4wjsXr8
rOjdwrlJ8RC2UjWqsHH2yn85rJkkA38KO064FQTZ9qlbaqJ5pYnf63N4YZUt8UoRgKU5O88PVfk/
byHMwpmQY7IWdbyV+fmTIpqenEqs9LEw6g7sy+uI2cIIdNqTSyI70jGLQwSGo5rKKy4oqLTHGM8y
wT7u2Bv+4lO7ls6PVDlSmWQRkWvClvktIBbW/y9NfUMtbc1uFOI7KOidRw24QjPChTcK9rYlsXvG
qV77olhp4Ss7iX069idVwYmMz0sApsAUVS4EA5vHAef6PxgFfkMgjjqD/hZIY4auz2SWrS7Whc/b
DEwAKa8sluuu2djPTjQ+7fVIJWlRxPryCou3IltocB+6cWtpookYx9/vx2C2bIqTIcz1V1Kk28uY
1Po7RlU6iW+lKcf92kEQ9tNlFxEG1R2L/Tsh57ZsGeeDtzQs5fhj0vnCPd1NiyYFz6jBpDsbPeDc
eNSw+t2xHY2zGCmYjqOMJePG7cN4yj7PcDXKG0zbu72w0E2zQnCL/sOakvU+Vb5+/099VBoCdJRP
h/3A0INh2n48elFJ40GWnS3i9ZpWYiIXflhCgc854lhJR490QMEEZnWt9SENOdQLkhxOUBRTagrR
oaf8hsO4qcTaB2WgLdO5fa/w6bvvi1CBOtc7uPCSZsRdmmEtPBn7vJGezTSnb71dbMbxYMlM4q1P
4g4lPzP0pBAm3Bv9wnHeTHbgOivtSjA3hPcv+iiaDwicz+44YsY6ZgOgXsl4FxaqjkCIBvgynaXb
ER24Qcet003cKJCTLQYRI7ETrNCl5s5A5ETPNF4CZcsbvVPs3kuO7OsD3Zl7MyzrxkE1xkvF09si
L/c2vcFjVn/XcXcMe5o3aJnN9EQ/72rG8dySXyqHD5Ojo+hTjGhJ0gHPAS9J5v/GDFTpPP9nEcdZ
39yP4naMZcvJFGryXMZ3t+7FOCruw98PbtaRnr9N8E/F1qESlL/qG13DH72TEnn9f6T+p+o6zBZJ
DcVwxWjFwh+U3Ci7baaEs8CseCQ+nuEBX13UeMvHfzG7e/dzMcqy5W7p9ATZxk/sfOiOGhfEdKCr
DEUvBNjn8TuejxGh9JM8gkc9wMIoXDqQ4xn1EfIPywuTtlBQDN5HmpoD1PA9zG/fWSkTGLr3C3g6
XxU3ITbdEiyvSjC2qLwm1P4nFLQt5YTJVH3S4NP88xFHovtuUtgKoNJI+PbsvxEw+Dtzk43zVwZ3
2bjD38Q+LJOg99NwSmu81APXECZc+uF7rerkNYrLOeFfvx4/uS9U7z7ftTB0xL+t4flkwxzYg8vd
FAWuEr3Nebz5l88ij61h+M/g7ThW8G7bkFgFJN3ggaWZVzBQJeShLFM1v3Wm0pBQx7fe52ELtRr0
OheCrl840RQFZExecW8Kd+hVntbAMSilPYqESnFVzMwDAzC19SJybElhBqytk2pvn2DnA8o9MQf2
ws77HAUV8i5OU35fdiywxJtoCciSST7Hz66bImVzfT6ifMkLN87ZklJCVMdqaP/ZGLlRDPn23xNj
kR5qy09qmJkp0179OSqpi9LkhOzhKZuyCvpWTmtdEGENUIH/1FmB8czaMsrGFZRJhuS+4r6QVt+F
uclg9IqOEtow0QPSOM+8prGbeQ9RJo2XJBdUCgCDzGXCt7sxnGiHBnAIccJaeUnngTB7ijC3xWcx
YtRqqwUybiNcZJF3QYWYmH3Utzi+WckjMYrrH7eh/FHvRjcWiy8Q1yMy+2LNhQWLeMbdloQfWLYH
EAZbhkiaqm68UGvOSPGmMI8gdn7XBCHiZTATaOpkjheKmfgOCGt8y8PABK9cUSniG8uaRA/bUXXn
o2Z6m6whh47jY7Nz55s9+mCs6v1u+MrdNrRJjxBgKqqwBHQE6LWtLkrhycNMyzyAhhTiEDGkTLNN
+gK0wvYShuErfyMVYTx5dnEKXuV3yMAvD46VcwlC7+7kt579U3G6zkC+PVbJEaw6c8NoJyq0CUxi
hXmk7whQAhhyTDfnyjrQwcX62iCGGt9ZLtpndC9CvFveyrmSTpavWDny4beoZ1HK+F4/9wBhZ9sC
aui9+8diPVm0PQSOU/B/KPT0pfwg7Cw7kFRkmBxN9aIxlNLEpauv7bR3CR/A/mLgjKn1jtj5yvRQ
FI3uc5QvEU5ZvhfoPhaes3tRTxaD+fUt1GpBkQgHW9WZ5Jg0YKAlTsLq5nntZiIOg54FyWvfPKa0
C8e71tg31Tqo3bU3uWZT82VF+bSkND7QlZBIphZU7eJiUogFkkFvHbCsBRcZ5ZVepNS5/WMPjKHy
KoVSYXx1RKeRKi/SW1lOrGdc0O8J0E7LgIiwNz1LfaqU8+3Q45EcTvA7FvSrLllXrSm6jMMnxqOF
YRcIiQw4wLfKSfFjMygJE9M/NmFii5YM/mDTFHWs5UlgsCkLES5AB5w5IX/iO6NPoLVo13FG4XpX
hrhny+4wRoi8Fa5kxifetJjqBPK3wN3fVm29ct7kplTQ6qrWt6wjI9aWmEUmDMLBzQwUCC3AjNaX
/gOv4hm10u/F8wdzsfq3KR5v99/35KT19WUxmhmIP9YhyALsiRRLxQCWgJuQq08SjzjiYNZUPmIt
WUvL3qzDLwKb5tBlUcferwW+qbr8bbgbFMmLh5Ckcdezl8ekcTo108wE7uYBerzGqXPdtkeshKtf
i2kihtk+3ByobCpHz4kJDuTQthuSFWDu2ZpWluYPOu16Dn4jy83m6r1jouCHFOOBw/6x2pTMVhUm
fynRLPvcivui8K33cO77Bk2Os66CWdk2eSUWcyWT0NSkmxQC9moolSjlNOLXllHqbsxrnguXf/Dh
lUj46LDfuvwX7rU53f6QmZ+fshF0qiO4uGq4rXSQCgX5bSJPhUAY5kZmCKJSkPhTN134RxZuXNCm
ljDXgTYbf+XDqTumztvENt2oZ1JjnSFwO7M53x7L24uSffT5sntXnX3S2pvShzTMHqvuv5eTIW42
hkiz3FlE8XJtNhDwBlFjAjrwswW4/Ee6FqnRVm4VHsFWgSViKq+JGmkgkptSG86Hk2cU7EfTj66r
Y5+W5uNXcb9Y9YoRKcyNzcYCS1GkfrZga2cf+/p9XQsyL9Cy3UoNy0E1QEm2OLdFn2XmFnY+Gocj
27PAiz5et8FnVFAEE5FjkWT0UnBrv7DmdPbnG7mNrxY5JE8lnRmCTkrqZWiWRUReyyQOPZoMY4dE
Ijj6Pv+UNd9AurpelTLD5tjPkWV5a47GRwTGqY8LcdgNXPkNvqb9KovU4s6gfI7NuaAfBW3t7Gwf
ZeW6VVpHHPTxfM7QIjeJUDcpwT5+sX27FQvKnlQ/o5uM1jOJlv/assscq+NaE/2IHfciJRVSZJ4E
NQB2V4UvNjoko39fdHy0q5dTF9Czv6d94V9fDxGpUtbMVZ9sEBtix0H0VXb64/yqFceKx9jZ3RG0
qqkUqvGhitPqLYL7jxfEamiF/JsY+ueJ6n90iFA8tSf7R4+1RKXsZtkywWyIFlz5VB8BEVLNiQrq
PtJk9+EgDPFWGivYXvTHmIaKUOSaUUjtNgZq/sb+GGeKM8Ct9UJ3Rpcurx0L7Ek7+cHNtl1AqP2G
QCuvKN+oR4/CJ/G5PRVdB74//ffektskXOAT+bLkbWFUJn/JDa6yqC9mJ4UAwTNV2cVKUjOA+twq
T0ZlTqqfvqwr+46/CeFIcdQ8dPyePT1+87iA14qBSzFC20LvEHpR8QjoOaCyc8NjP1T6PL3Y5sS2
Qa4H66qqca7SjfHPz6zWVS+t8hjSaDErhoeZeUEgDFQuMPaDs0GVzv0EtX28Nckq2AD6uZ+q60jE
ztyEDcHMA+JCbrUhPeJx8p3QYrkkNKZQ3Y/qaUt1RrlNkRPNP5eMqU5nrCRKovNUqK/KQnLOuNY/
6BFfm6KljiNN5bxsIzEWKIguPPVJbUxSlXTSVDiIUIgk8nFaNHQQqTBAyNm80338vNuE0tO9OgyM
xwLySQ0N/1cvhSrlXXu/4CnomTAlGtNVBWT4bOVlQIkB1dSlSUWixFMDhDtlMH9sP88QZ/eb9y/Y
E86BGVkUIbiJc4CeLuyfXQ1iTVctFkdWJs1fgBwb2mRwuifd16BF2DJu4qWIT9XSRBQMni/TV1cn
tbDLQDoFvVbZKSsz7MBfApO0/blMcMnR2FOqQDHoTBLhsze9gk+UU7FqhULj1fNcTmB4GQE9q0l5
dqkwSU/9gaIdNSQYQiOBqaN/EmLsE3HKAcsyoSLxaBmGVL3DSBPMrODPSuX8Z0P/VxMpKWgxyXGc
/T+Rz0l+64xo37Ws1fOxKsAS9YwVF9NuPr3GtRH4ck2ZVbAzy+jWgBuFUb1BiydEdGOfRmVsnao6
YhlMbN9ZWNyCpsDcQCLir6DzWLvjN9WXXq9pbBmcy6e3EgPJEgfVRf/tT1D3TIvK/kgrhc7Kqyou
8awdNaPkbrLPgj7iTw5plmJhS5gH/FVMqY6nJ0J3WeHGOIWMUR64+gQR3TuaCX7rg70h0Z5P/7Yj
W1kLDv57EmOrqpvwFUvWyUVHq1CDHkYOfJrw+bGRiDW9dXfgb4AF3okU3mYBAby0q5o62c5/jWjN
sjT8EfILn6GunH4Ae7uPwO5ndbgjqumI2jAUTVo/5vbVA7Kf/eKgCM/7CA+9lZjfaRcT5GncM5aI
3GnqqlJ9NsWrcDlUFkZgF9mfzTLZZ9xcyaM4rubb/NbTIJ3H5lpkfiQX8FZVJqqnzutBDN/bwMyU
CgpHnGLuvMmIoNWMNBaR2x1Gzaofr1NMVxQouUilyOO8o1OfwtiLSCHE/GcWFM6iPBJIc+zXPhqT
8E2BObbtdx8asNVB5JMgm2UJQrcGS8PkKCIoPoEMck+au43roTydZKnqSzqgxhbpOGrMFdA3QKNE
mz0sc0Cso5Iso0Rw8EJpUJf/5TuECVx0KvqOMkPQnaUgGyrC9tUs/16qHw7lvK1UVI1wVHU1Mv/q
7G5q6QEPich2g9/LOjoqTpD2Esr61QUWsrlvkrAlvYSsL9Vkeo/6F71/reMEvuHkkckmnqCfN8RE
+9KHpH3c+sEgOYs6AkO7okUyg3xIb4RCZaLO3LPXerkaZqnnBDrxb0QQPLKRXELA3Anb/Xnemklv
SBH995gL51uuRCBUmbwUd3qmByzHv7qeDDK3vz/m7u30xLEqPRV/mLZntCCKMVc3cbGgFZLSJXgA
xYloVmKb7uGRlKHvnI4q9z1qNzTA0y7mvT7lHxPxJQtifi6xKwR1oX3j/DBtadWUfXcktvhVdlY1
3V8p4KroVqAHzpSGTySLxaai2bzjT0GdDS0BV2TJn/rSsvBQHPV9fruvOdg9xh5VsVKJG7jOkhp1
Uu76o/orOdyNj0SxRmjGpKtmhTCZpX0n8w8cvcHCN/lzaZ7xrPVx0FAAgWmElE0+clBMLnNk7FCx
AKIOZtlk9Peeqq72FhfjLfih+Htse6IZSpR+P2cEJmHKc9PZINbzhpoApAPFlpQHOOFD+1uGM+pA
9bOZlvCpjK/tdvjoZ8sAavMoRV92NUbXcKLnGv5r3R/RTyUSpiHzzJVYQwQoEEl7wAyjSoRzOw8k
Lh98RrD/os1pN2gwmuc3vGXbmozaMDaz4rWQjTxa7NkjB1uxFC8QMGMH5bCqR6UCfSRfDTEsJkdY
gencAgMpzYlANSqy2uBDiPEG6edF6lYY6rnoe5LJLbe3iiUgRkfaBUmNitbWJibF6ECK0o3on3nH
bJSaLqhGhC684x5TuzKtIQfQK1CUM39OkVgDpinQ3E85fFHo7lABKIcN9QEfeod2EW6pqJW+QlzL
NoceW97c7sEA8At1IJQS+c4ldzFc7n7QLVj4GtCRWFOR9lmqfWSpbVXle0x9vzKt8TGOGJDhRBRk
V/MNX2foAHYK5TBNLppHyc7iNAMz/LVS1Er/7Hy05R3vOnAJ6UCiCoOYcP4lBGnTKAEvmX9nSzRd
soXVeW+EX6yt+cjVzB2eFD5l6dbg6CjnhPTj+QePg07iYIpGhQeEVVZmOio4vBqKoVJq5OwR8zY+
M9GVN++M1Jg1aA3ly66cD22rMXDBJZtAjROhh94pUECzT5UaVwSfUZj2JVr/f3t+KIDtgms+cz4y
Q4khRWWZ9wM+axjAynwAnlSxA+gWKPcuSc94/SW5DLGz9j8sabOLvBG1grjwuWEmpAZrrf92A45U
ZyFvn0dxo8ABDaAiOyKNL77x1iVJv19XdfKXTB1rEGBiJr3V7Rz8JBiD2TwnqiQ7GFnJUTTM95IJ
i1iJBnLbKA3NiPVRNwbrAPPfhUxYos0tBLfrhmAodKxt09vBMs+iphh9R9oUZuWKonb5jSXN14ia
zQ5rhRWFzzJvTY7GGF/OMD6b86leaWhdItVxaLYn5GqMEfOKeW5Y1PWRkSSUv0p1fjb0+VqcH2lW
qF9V5KRATGR/E80jwjW30u1UQjhoj7imRJ4DT6+BUoQT0ivfq+9Ttqal2SSWU0QY4HaIcySMFUGL
926elayuAznklO4U0H1FJqlCuSnirFnxXVLiw7rARzrL/4OMULDBWo7PYYfmCR4S8v6PMKOnsixa
iKa5FNsnTwxDUtmMTAMAsqneeE01QmXAQLnsCAic85QtQTFeyEr7eS52Yddkn9Ctl76xeCoqI2tx
ghTids+xqOj1PnYjf2pMk5Kc/i+UGau3LMWkUNNXmNkovVyxAVAs26x1r3T60/07VCxcnJzT1CQ8
fLiachRm/WiQENpswPQE3UYImBdtpBG37JqYtJhONzebJzrILylI3VJH6AKKIoTqZxbMOhrD+utS
1no/LngT1fQq/DVga8VlfD2nB/LK4HRg+EIwcb4T9z7UQR70ggeS0nqwcDpLEWGG6ZfuyC9N0RtJ
qwpi7QCtJbocrHUBtFrUmpel6GrUsvEf48KQTtwqn3//htIxGmOLvuKOwu9x/2pXXs51dm4gN9cZ
nLqsL/aw5oApScCxzKE3zEzDw6A9ZJDk6b5iy+zgSpyuFYIzpCJf6JdUVXgaPLe1LBykaYeiQkWS
RyzuST865qoazl6ZWncH7fdw43gSz1sGPswiwYW30JUQcKpW73Apu6UWctBCGBGoxq2BbhAB4MzN
NrSmD+ubA0ZIRmNJT9H5aQmvQmmjBAstuBa+m//k8/Lk3TDDU6apTrH7y9uZJ8we+wkvuPSzrpcW
X7OcVm6TPb/8ANgGeKXYmpZR0RsgrCcx5GkIu4HNUuFMvEG2C5GdBC98ggcI6tPtxHAaVbG6125E
RXrSlsC3dT/1F6j08q5UxkrLY43byscECAiLa60KGVY/ZHsXNOatLruRBNFOyaMgAdkeGKBcWEzJ
oAdn+aNEC2FZYAWMknkdcYSM5S6isOStpsnME/K/gkFxeLfvOFIyITgdXWY9LIOpT/niM0+L7Y6Y
RN+6T2gDRXVhytle7QSAZdkAqXBv/PVmqvG1vnAeGRiQWsW31YSw5ZOl52Ft5Zjt6JrWbDJyEK8R
xjzPLO5cJW6wWbDirChCQEdkdFkeZfUQDHvoofdHJ24QvVGvNQpM6rxwonf+JAeWLtklacN4M7Sp
0ffj88TEihFiKDwsLMVxOsHNbxrr3Ay+HMw6GYNuWeRIDjLeuf78yyALMDHNg4QDNeAIXCXensmP
F6Vi+GDElma3Qf3ZSXI1MufS/LmYOdqrMs4TunkLE8iJenBALIFCTow1/S7BD5z9/0IKk6QLuCsd
ieNA7A4iCqLx2PhrG80xkYho3E/Nc9roK1DPVl1nIPGLsnxNSK1GdvkmJdlLqBC7xWB4KWfIY1Xk
lcqPi/o/jtJd62WQV44yoo3dApN7bFXc+kCZDb87649gaRJ3fOHKi2c1kicfmz2AgYAhJ7mcEflA
PH7sGEEf/zyT7YiILtHlFfYVcmf4Hiqn7y4A7WWeC0zDX4hTX18/72vzbjf9dzoTR1UHIxjXdcSc
yJkQtXfbcPqAElEz9q5ylgfGK2VXdyxT2J6/F6FCCrR8vVD4vx7dRYYQcRKgMz+z4YcFye+4WIBj
TWfx2wGbML3nhseFFtcDHSaAzsS3IB68eAS5603tGGdUoj5uCeL7AyTbIJ5zzuF6UvRF3Y5njNeR
Bbi1suYpCwxhEJBjiqaXglocPjyBr7zXjTvZfnPXmTC+ttG18WYaETyTp62EhjpOAey8c8K8ZKXm
h6q3M3LMWcPemz5J0kNP+fe+pBXD6bz+n+zx0huxvvKtI1WbqxNkb5COflKBoyy9xdty5XkWvFnV
8K8I765hYs13ACu57eIpzJNe546uY6211nzLG9otyPTcxAH/cOI1KV90se8PVxweVSythIiwFLe/
bUi9HlHxT+sgzTF/u8DA0kOGkYmgLKf5nm7+fmnVE2zwqRVUa0u9j0MjetT48RLgVquHe5lMbJrK
TJ32ImpjqfvuD7cehzEaBb206npoLzpyadYxHAWdtueErfmjaXX+bwtL8g+ZxibGHXpvInq9Zhqx
s/g3LmAkjnwcPhYbndhBINw2Rle59s4/KN1hvktgDhu15tRnCQLij6Q5DAUvcCgLjZJJutq30i+d
OpQy6xDFc4/+OfnWwq3Ty2t0S3M9wldro5iL+mOuA0J8s8yUi0+65xPv4wZWTlHOySio8PtJr3t9
91IgEWXfNvmH2B1wuskDD0mqw7T3RDY226vzeY31dM9qVus8TRwaMNHZPIFCiyxjuxroPFk7Jyzb
r0uVDVjkUKqd04cRAzTkfIBQcSdl098ykVHZK85t7SLX5TQFqsGExDwdqFRwlSZVhFXwhWcCo/tt
guE8ku54fCD4O1Qw/012xziXjgblMyPxW/GO/QNyUEVBWZv0RguPanbwtoNC9M/Lm07E9oziXOHB
rjEgfeNJqs1jUHhnOz4v8Yd4vZzwPeFRs9PuU3h7qkCleat/r0SOR0su5cZKm9zqG38Mx6bPUy/s
NPGDE8anrH+9WAqA33uJqv3t92wzwaPWvzOLfXGibqr6QlX82gFqNax2OVqtY1GuH2M3ZwQiamhd
oQJuAJYmkSCAKp+z/SVsaXVTABmHdBEHPxK7Kc8gID+XTFb5PgGsu/wZGkOe434B7uU56/iTRfwT
oFZrvus1+F8G9UdbyTJsqP8LTbiGjhU48iX/q5g5rpJNnH2zY+bfmvdm/YmStYfQSFnKWkP9eY2a
B7tV1qetS0gg2gaArrmTlvdlVxA/UNA9ZoW1r9QFR+aE7wKa8k3uqsCL4KyS477gq49RRmVikOvE
tgTnXNhqmSe0szoDSo6baI/6Yawc8uRFeErB2GOrMS06a+uWR3QnjrU4mYVEmhrlQkwNLdyohjor
ic9FdefrfLNyiCBZBTGNCtlRTCDlVChsYQZ0NfC+p9qxh0TsTzIf1YLAvbgEWQOnaOieuDVTr0Oh
b3llc5fY4CAL8eNV5x9ElP1XLPR26TzmbtQy5xQwivskW7TeH9HanijPNmIxknCqvzzd2ihpBIHR
Kxdy3q7daPOQXr25p0sVnwoJCTcOPev/T2VJzNZAzJP7SVMt8ATd4SR0S8IoWnSZsj+guWDnnQ4u
N0vuzbB+eJNiNxXQwvbzpnJAbUo4eojFOkw75Ov1w45kNG/SHrR/rYdg0z9aBHwfuN/omyRvCSnK
n8NOuhlhMtxcXkWWnMS0rBXlRR7NmU2OB3PIKFES3RVX/zsOUzOsWuZGwrkUd6Ep3XTHrn2OzjFz
QEZEHsvBAfvyfEhgg17TN5vhHTYsO+o0+vNp3TPiI2OFcH3ySZRKcoPdGS0zCKnECNHDYI4YTE+d
OUalhk2DZvCBluLRqZCtcG4k2wHjD3+C4xnAjvq75AfKQth5AfwwSjKVEF6YlAapDldxbekrU5oi
AuwS9QciVXViIdHfqft+OH1eydZ+zuGZPofDCktMrh5kNcSWmgjtetS2Qm9FGTzvC5yo3/GilKXp
a9yerI/vdsfI4Kj04wdHT5lnEpwtQntmt8qiro435JcDSPtzHGiZ6jXy3heBi3UvmjRXXTFySKVg
h+J04OI6fdtMjwpmGuutuwvn3Ga0IOJ7nQFSiv+p20PDhefsRIHd/qXzdl36RULy5fpQ8oHw5G/U
cBzuLj0YLq2qXTbjluepU/WYD680k8TfHknCCvvtJaYhxuHsmkGiXnDf7Ed4WAJuV362ZiO0oSiI
xwkc2gcJI9VgovY73KUpq1pkFtCl4BQ25aIMTtb6M6xveUxLjnTc0nWCJzY0KSZqWtz5NBHNGLNp
s7NC/XVT4OXCmkINuyhgBFPhClnsp9gUYmF1dpO7bW76sFsmOqsITG2uCcGH9H5z4YW5ubO25PlD
rNGsuUkxxw9ckHdKZO+IRDq7dzb3YwDcNw4/VIe68i7I5Q8E8/5B/UP9MFd+/PQtJwYOI59/gwHc
pCXDTAbnUWEzaDFLlX6CReRbrbbfMY72GdYBBhyDiwFUdJUP1XcHoaeVoWB6LwBssrGthppkJLGm
M4l+CsdhTzUVJuS8Ts+BWa15JyWk21VVKZChtz78BmIJva2e2sqktLig8ClTtFBVUNfH4caX4z8T
MY+JZna41TxXmIertVaeHhqWJ0OiTjVHlqpqvq4dGwxMZHWsv57aJtNvO3Q2P419IEMlXudUz8xP
NgBC1pJNepbOUXSDiR7zsgTbj4KvdWbOQL5fd8KTBcu5QYxlTFq7GU2luLpbDlgpEhQ/k09nShP0
DNhQxqc3XlGgGWTKqpAbOTthsU2+c1oYjDbSV1bZao7rbNdj7iglwmR1OsDjMYp9l9jK6y5UjqTr
4ZTg0cCLvaX/NsceNBVLuqhWyJcnPLrHnQ0IVjxbJEBLP6JLhreMGUalicQzh9Gegw38ZLZqsLPz
uZvyfyIHRqBoCziNMDNffNalj21e/ZyZzu0j0uF4+BsYw546M4VAhWqli1S3w9Q7CJgeYIP4R5mP
XAgiJPnTDJexA1BNvZ2sbjPqxTovUpSckJZDFae0ocGTcWn1SssWukoXXjoqR+EBCJ64Z0Wb9Q9S
t7YLkrf4cSKXC+Y20aPRvVBjGNDzr+6M3FL6OwU1SqEuoc0ny1N+GCNVYuQOmFwUEltThEs+EqXR
0DGoyxux4u6hgTdh4ooz1JEhWHKicH2wkq3BqnSbQeoKx1r72baD3F4CBjYm/4CKRfh/AR8WCxYw
AfJAtGgIAa9TXOuINGpHlIpu9DamTOnNTcuLj+QN1Gv+kykZcMHG233U2RwWRk+JOLPMIPtd0NiM
z8vV41wFutm0O3Z7fTJx3CycQVbthFw/AwiRdgEwi1Asw0f3vJDjHVfkyPFgg+xWQBcvDKQOJ/t0
ckmy6XzL34O7smUbcMNKFn0/U98q+dR74xtBj+kN6PpbWM7ujkPNWQJVInRviPULnaDiKMif5Ol/
+eVhe1A1x8BKxmDEOOFV+dcGKvuclwKmk34YZrQufiH9wBuBXL6ZJ8BemQd51XLAUyokO5+u7nKT
eXPMkvWm0e37DNdBZvJXR93QftYxQJ6pY7ca0EFOkyEwaoV15IQWEY3TLS0EWpox/lW8n+9o0+bk
GaCcRPHsHaXzc9ZXc8yhzhIFZJhRFvym/ZW+isxp2Me3BMhM3eEhg+N8u7WfLjbacrBgYN+HBwKd
g8pdltQlqOC6sUogWL2YSE6j71flvGH/qV9ai2YeCPi/to4lV6YdAkk2m2QlZ7RMLs4Ks640Qqh8
6wYxOKaCiGo33/egD+n+tuucbcmxPk2680zxvKMrIh4i04RfpUZ7G/JxagpxA37eq96fUwka/8kL
abC1xK6pl5Y62eF4zd7PPMrBjaSNSsT7kHd6cI/BFiFb2cHXmU3PuKguIWOSH20tyZEMSkUtM4PD
dyNUVgNBS8DDGhWFn9fV8Ws8OOR2TYMMkMIP0ua+qFtlBlF7P9W+7bXEQmeM1fqzIygQBbwDOEGh
GJJaErvXNucircdkp6Iz8Otw6ozqlxBJQrvKgsKhqcQ/6LHgULLF/u39Rj7iBQuXLVAZWNftRX1g
82c8ytf2IltfHvfpu3tQbY1HY+t4WtunGJAH0ceoSL/vCEX55GjhVZS7+y44gzyO4geZpMUUZi6W
lZEgoDyNuAG4VzAn8qDFF8D2Kc5zXDe9bZDENCHYyNtYxLtg89nm8t3wjt0SALJND6UYkng/WjpO
UNP4QH4dS+Atht7mdSHRAId0B7GYZnj1Tlmi7ObODclAgTa1GBwnZhIcS4cT/kzdK6Q2xnluIC1E
fn2VFw4Zd9FYzrbk4qS1avZN1Rs33f3nXpuVN3sWv5E/khEXq2ybNii3kTeX3mIJB7W1DWF1PI3Y
DHQf+Hzodf9zGC1u9DkPtsdL1stcgz6C9HMal53oKvtuz0BzPMAXynj6m1Zt4tG3D/MDSWq3in4p
fGSmPgq2kCwbPQeJewjVco79IUeURcBQ8Eo/5XyGA6/l6c+026j/SfGLIkq4VZ2QNWWnK1AE8viK
jc+/JYRysTyx12nwzrQXVkaxxHCw2+vfJ5llk4EeOmJTM6coodOXc78wyyJvVb8ZNLGGcsz3uX0J
6UKcv583JswyooWkK2CSSffcRjsGVDkFrxUC0h6h9x8LMLsOfprCbj52yL4O2Pn/2TbNaScCzpRk
eeLz1eiltoq8tRXThIskQarfIgNuwShWPN9pSGA13odwI559jn2GT5L+apFaQvvlIAlvYva4txmY
aQI30YzI2mo8cYJ8DutaM8DbjckKvO9bhHwAkFiDg18YmlStp6ZYVRYRmlyjihpyESyLK+xcO4Qo
oYyeXmteLiJW/z0RZJ6ZFDBOS3fnb/rUjrTH3Aw6XloMi4NkqQb7p7VIswaCt+XFUgZdazb1Hy2M
MlxtoBZOU3KLryxw+DdMHH4F1UMWP6eq4aPc/mquo2ibX72URtkCzKrr27hIx3gBxCsMgkUv+HlU
mzLcnm/z8C4/PJLW1xx2CcAzAdX99MH5qg5Lzd1XubRFSKadRTXtasUr4N8+Eqm538fzZ+bO1lIp
8CdNn1C1szKs/GoCr4m/rbJcGaVw1mXv+r+TLcELULAzC+dhhfai+EItikoxMCy6P8/roZE4D4NW
PMOMMp8rPfj2bjWPA8rLhVZ/kleHTxWSgubQDVQyj0A25r1LF0WCH98qBHl5vLA2tF5inW3Spk9+
DUfqBtpikXqMiLdKlh9wuVuRK7RUqv+h5pF5d9RgePMOpYDaDg9jTNxOAK18Y1ygRtTDqI4x5pp5
/APshJvTz9Zb7pIyTMacOvlS0QcqeT6ajJp1Ys35R7AQNdH2ReJaeCPvJtlveQItrmFSTRuW8cj0
iX4HOOxO8fUS84Eb7BQH8BYKuOgGAJP20QOIWErAEWCb8mlS3VbKaNgYf0B4AKCviicMsuQGLcN0
Z5tsB5msruQmlvaHr4PJxq68XATIwGFkcj5bAPmG06sy6TmnkbF6ezg6UpERsIDz0wmzspLZLXcr
r5iGHmRxfLqNuKqM3eBsJ+5ADP6nYSbuCCFWAfCTeJCVWkONU1Ljd5l9ph6pKfCCl355itqg+OWX
PuoA9ZlKEwo22APFnLjQEeQ8ljrZ7yySTCo+eQx/b/SntIpuQxogwZIOuHoQgCVaGryLPlNHKaIM
xhBlab7MtpRsm/0pHzAg8suqIZs8YTBHEyMqgv99H7nyA0Qzyccwz6yy6btC8ITiKeisz4qer6wg
BpW6R/OIaZzs4pU1+p0ZJ+FidAnVgnuACVPWq0c0iEoHtwcveVWxcCYl6WNDFWbVvSZ1fI8qP5c7
Vm7+15eOPaPZxcaA72crTP5/ZrhTflhFgTWMpl0IwQ1d5AhQuObB6rXDnG/nb6e5eJkBvLNBabYr
/bxxTjp0Q8cIc+06PYYPoKU4LbiQTNwPbP1k8U9M42akvpL2nBvi7XCbHnM+zXEedPAl0b545IQB
j0qJoTG6uJKN6RMCaTa2qAQhd75exryhFC13Ot7HFQL8OGsHzLgy0hdhjavf1B4+1pC85zL2l4t1
1dwwnn/CWwsKs/R8TQfRq9RG/wVQtiMSdGW1P7cl0jvGa8GDXSCKfBOvFwj5zOC50IVNSettzI2S
tCyY0MmXJapz+YkCroVoZiu/KUqlVBXukRMGaDQdWkjJSr085EpfKA45emKR1vr95340bIQXcisH
XnagZKntsZVS0/Xv3nvzg4YjV96xZrxZPQbmA0+8nIkbuJZHzGRSx2JjSW/ZOoXjGXYrpqB7yC/Y
h+fr8nTphVz1DSgs814VH2XbtIrOC/5/yM5dtgL92Jwb01AKbt42Q0PzFP5I6esORcolU2NMEeMi
m/CNO3Pu58Ew5BpjrgHYb0x9h0ILddnstRHS9u4tM84HjbgV1YoqH3e0D7i8L5JhuIJq/KBMPS1L
J22It1DijLj/XWcXzQIVEmBvIQ03GiZOnI8hU64oPsAs9j5e0NDZ3CAZZiELma2/+quene65vu45
vgQEsWdoomHVSjHF7tanKRvbKdNMGIzru4CeyEnt0VoZeZtXCy71LTWbo16oa4SLNu2qKZ9w9Trm
FenSAGUIdQBMlfhrzqNZpgp/Vj24aq8ICr11I1pxvLPz4y9PoUHMqUemq3xNfKljwbzfVAFi5JQC
b2T80QpXq5dVks4PcGyYOgT8FzQ6MTdn/O0IxLSgNl6nFvRlmNoSXRBLmSlcK2VJ+bPa95VJqNqD
pVWI20ZRvMZMdRdVKOEfSn5M34MFPxs9Y/I6Kp4Z0XtF5OINR0f8pz7roMHR6oQbR1c2W2CEb2YE
6gW9q2eufvpoAAGzQ5Kapezb+3eEq2gIA0EzRvpWZ1NEn00k/pQ3tbOpTn5PvNw6R1ilBi2DILa8
1c7Y1E3sNrig5Ke4bL+yMabtKumNhOczzK/kubzpOOzc5O8Hb2hSzgAXwzKYUm8T2kQTKcG8yNhF
Fm2D5qnXloGbaEcU1BnAaFzBbVKA4ApHlejHLDpAoME8NPUtvo41KvgB1Lg0DDCWsHW5cDKd5LCp
7/h7PjK1NPU9DimiBB42bsb+3aravr/mh2k2FPi6ybPzvgrlaJU3R+9SmvzsxlQ/A8DC1Tg7atbC
kJ99Y/OV0CqsqZ+DORfEhCK5zZCTkY2MeqIxm9qTqACWzguxIejMLGJiAW1yA1CssyNhCgF5qRIY
o3IuKa0uCvgaZGFIhpGTxbYxiuboNl0dHa5vLTGQ8OlxB2zTeKRwqxhEpLhtLfgKzHAcfdGpCLUo
zkFKthBMlu/5jnsPW3/4h/M8te78zWcR1k0gYhsQJIFORo6iSuCTfZfERdDMOOyq0SxT9+vLn++e
oyrh6wJe5v9jj8IP/6OroSjK2VnjvR5YG1xe2YvhwRZ0jyXFuS4Dd2dJrzPo8kJVatIOt7v/sWXj
1WqbX8ehS+8liy/sdtox+cjFI/JQn7AvoNZ/a8Uj1HRMbjKxbtxwueX12HSjLKqClB4slMgLO4cO
rGt49XDoiUcbIMWa+w+w1Jz8Ctsp3pnkytGT+lLtd7i4E+PV1RVcca+MN59LcVkHhO9zOecHqYEr
4ypqRPujXvZHQ5BgzzJ99aFSML8/17BhU4QZ3/a8LWO9yAWmKD/MIncSmeqzj1DhEjH5KU06SFyy
gFTp2/xin+pofgNn9LOQIk4co5CFHSlz6luL7v5hiwGAxj2pzT7Rm3lQ64eHb9E5oev7eaz3Gs2M
x9hofBdOxKXJtPDJWzJuSjrjl4v2sQ3Lnok8iFV8L3O/x+GcsYEArHkdoBHb04ciY6/SATmvt46I
/FK0QHNAtlWx5wSC+aH5+qUoi9PN5Gef6+qutQli75T7VItzRjaxCy2ZBxpthDoWm5vMBV527zYp
ib3XHVVO9XCFIKdpUzgE3YXe5LD1BdKDGin4/mFmks5Llrm9QRPTI3ZqFMFObslqhZKmz59ke2Ho
xHSnbZOH/L3d5YabjyyhD1lhhQzNDGugnZSTrLVcK5wye6He4yUPiRBJpT0dBQXW6MojYZRF9A2a
28xCu3lhH+CLnAR+3FqFNtFW23MgVh5P0W7qw80Wvw0kg/dqREdfm7v72m66STJm+mhrjuIS/2Kd
tYj4UA0rGjGhjAaQLSQeM8r+HZ1KbP7qlwRwJO5o7d5diCk3eC+xFCFPhoMYCEvXHi5ADlrlAmdc
9Pd2f88EfSv4FtiyxH2VKQo/TnDTciUfyJ6LOHg5DkKC19l3cNDW4rr/A34QTLjAW/RXHxN6PlrM
Zpi/ZSedG2+NP9oADlwOSxWrcfrOm8STVJWUmJ58u8qH3niuwI3elatpqYszTsOS6ih177qr6NzY
vWl7diYDICbVyFJQ4B71+VR7j0qbrlwLRzyFRQx8yv2j7kOnL74DpuJ23vk8LRS8lJ0McdaO/U/f
EG1rswotbXatn76L729FjByKH8IyOeheLk5XOegLqzlYobElRfrQhcv6H5fAvIMbMvjM0VoUmLcS
WuQisSHXW6WBy0V2TFhdVKG3ZyMwMCEpeSFBmGN289o9YCD6udBvpNIsmmuoABb32HiqHOlv2zBY
DCdi7Rj2aA6n0LX6wTLRGYsH6kyzFXzIDpcndGG2vIHJuWd11PCJCGSt6Mmv4AOg49+hBrm8NdlY
WP6d5uAXhvk8berBurq3Xcz2IelnXccwtN7V3KBafGJKiZJTsJOFtjw9oaYfvYMRPNEP8pBt2MWq
GFWXCdREc00Ds0WdcDAreaUypyFn5zWiXPcoaFPVTI8k3h3cMvElvwCCzLqbsK4DOVkd9bjQEJiS
LP0W8bOyw6BAQnrGcNTMcoMtQjZ+MZJQSjLPX8tSnINloHRrsOOCwI2na+S1EhQazWHrPTkeMK4U
K5wirRIIBMECchpol2H/6htQPKS95OrE9Jh/ilAhYKF1kbjcA5c05EMLV5uwmaDx8czpbmRg30Zr
YnLcJkBw/GNhDy5/uYPSpGkKZFOp3Sbmq/8ZTRTYa+h1heladTStMmmF3GP1RGo9TlOTlSFIYm8G
GNFMu1cvwaVsHCn2gOAjPOlAzEdaG1fJkF31kv+517Zw2HDIsR7q3cwIJQSFHQkiWxxOgd/LNDoI
U+eZ/4AR72rSuH1zXcRulboUjzynD9GpdrgP7FezoGT+W5jQD65gDRuLmrf8kJpcm1v2Qlhbyq2y
OBYl7v9sur3iNffVNH5xXR3qfQnOENWR9ZlLIsEmIiLmGdYLEIDGBVDzkuMd44IT/6DIczNnQhcC
HcIeqZmA+NfWm7IoMJSf2RR0/rJrMQTiMsUjZT5I7Bpy5OQAx5Bb6r7jDxEDBhox4oZo8zgrShYe
F+yqJ/CZL5TeDq7WqXaDzgB6OtFMcqF7TXlCKQifUfn/OF6TCi48KLrBFr/FbEMONUUE985CpcVi
AbZdlS9mknfwpNFWYq9L0DWGW2Q+8Cbh9Rifp9zB+3J4HgY2VAd02YcFEdTwLyTvDgD7XCDQlywR
AMnSxk8iy1pNSyqeb7MVXmFpvARb6k21479PGs63Jxf3dsVixMXFPamFNN8Fv7oqe0yrnsve/CQk
CJRRygfoLNUbwXMuL/YpoGVJ8Bd7l02+GojiGpIL7Aw/rKbK1l3w5ZEHt2Jndn1uF5IRIWxD6idM
u4h1Rxka45+J3211Nq4l3+txCWvefnyIq/zzarEOY9MW1ZSlBfQPzWqUGKrvrWM/9KM4MYfZPe4k
yL4V5pKU8a8r0Ca7dmkLYok6BvAVNsQ9deGyjezZTw+9eyJWeOmzX4NgIdRoUQH/UuH9Zw5r7cAW
/A2dBdx9hnrADDEgDBPv8aulTGEfueEVb7ZVlW3kxdIjZu7LXnoU+nVFImTpiNRABq0KcqdD6Ny0
ieQusZgkKCHfPam45A/Ic3u8kRFBLVeD8R8mJFe2fdhlYIW/Y3yVXktHG/4PVe/NtBs3y8D3yobz
zsqpENw9gOsGtP0WgzJY7mmPUYc8oUKcRYiTud6grymAkw7EedBcEjDc3/4cJWnwS1JKxdh86cbe
TB7pscn5ZCFFA7/txCtBV6mI8TXjCCNYg+dZPYD8ScjZMBdhIrXAn64xSR4iRoPj1BZJQCJ3Vje5
g1xu/kgNAi9/lfq4Lj/s1HTRHg7sLtTP9ewGU0B7Ix0Bm2YenzxW9+akasS3GSr1WKpwni3RjgOz
YZfZrUlkLR6l6r1M8yyNSQN+s/ZtJ0MTyOzs7xJNquQsUhEVPuPSTYFEancYHEd8hoqD1+UL1nAT
Kqfl29UN3rn00u5QbZbUES67V6VTTrHKoKbVQbU77nTTD2Tohq3seldikDwINkNQE1CqjQtwBj+g
graAnhA9DXVEn+Loev0c/bAb7+X5oZkFNvTq9bMOQC6gMeGDDJB6/4WwltkYoJFE91GXFBnSUpSU
oKusr57d14cS5S6XyZHvCy+SAZqPT7JsKcmyfcKpO6RvbicBsM+7+4JOwyTf6qkbVNF3anw+3J3y
UyVWhLqewzgPlKblsPWqgjhGGWHMZ0dtkUdgJ/nhmr6wZSe6RqAf2P9Dlbe1I6xFfDT+KP9rrXpO
NBY3RTixuFSs/szCrJyDrFo9riV3uRsppW4oLk0GZXBUsyYuz9igICfoK3OnM/uTtWZFY1i47vDU
YDQeCDRboE+iXlPCehKCngYq7vEZv7AsXH+ySyIXn89xOdps83HzwuAOok7SF/45/qLt45N4DN2K
d9Ouh3TPW+N4iEZlXUOMUlc29oF8qrMTrB1oJZBzuGPl8MEQthKvwIahNxzM/10O0YT3dWLcTl0H
6DGryGCyf6TwIB/TqNYZRfT8oaA4aG72Ybouchq03Sh7Kg9NA3nOidr3qZuKjv7yvFAGaR3jq0GP
3GUAVOjRuCTYB2bb4hJ2j00avUKyeLWWlfQduQd1rhA3pCeSf3vzbFPfvZbIw7ySy2ittrmhxzvG
uuro7y37zZoQYy8TO9x1qhU2+cxu0DEcBBotBGYnX3UHQXd4c2MCS+Mg2CgIe2W7SQwrCOL8gcD/
tZmI/Gbf2m868pPudbkPPtT1EntHLy9n3XxlIgRL0F0hLjk/ke3e1uVxf1uf6e8eNKgOWt+zYu2O
CEhvfcaoZgyupwiClBBvH5xMD5R+AMCbrWkCXM/l4G4rhI9RBTRke6nOlfbrV4e60BiModEdjFZq
D9SdbPf6ktUkQk7lEinkk0kZnxOYGFnq0vwKykQS+s1WWacNKkHhs6PnbXtWg786iMTVQw1414Ke
K9C12mwAiXhuQzNMnylmAR+1jgVV8enbRtvm05jRSeca7NIAFrQDfjyhWoOSPbVXBqKCfb7uM4Vl
/eyq6MrKsVGFUuGHN6O/klyK3WDVxLBghzvYU/TAeIVuqWBh8ul2vz20NYDhAZ1k9cILsm/wbJ3e
cuoquqyAFQLP3ulVrI9d2x+8LGTtymI9tF+3Te5lgx4WlsHcI3rJszhn6IGOqZ6gt4P/79Qmx9Ki
hZjlIgO0nfUEp8ec5gpRzuPXcgf+zzEteB1q+PcqRwpN1yk1V0+AOZGCtBxiHsVvhunYAlC+5tHW
ENmx78wvATgN691wldX18PXFjwaxusSRuhIwYF8drtYyA6m+8z0N0VArFPVg09MTEzdYoVPlMAdu
pHFmsMPDwz/IR7N6EHq5HfJ29vGMkXOnB+9DxNDa9m8ggqdI9OmpGdCCl4lhZKALJGrW/X0mzN62
0qsAgx+b3efgvN3mbkUbjKYCxb+EedH7vqCPcBbvSzhf8cypp5HYG2DJuVmp+H+uJehcopsYqtHW
DDr68HU52mLWIBmytEXmsuFNaYA9xBAjrEPBiCtvvVHU/b/oSVu/VPkDT+K+jwrw+Wq0/PIEsSPZ
OBS9NMYVVm0w3lWRYSwOGZKlO7Lnx4WUMYEH65rQCOqwWxIeScLotD/Vg/wPjRzMw508UNDQv9Lw
cpNCKmqH7q9lpTJltWGmVH+blUlGQKx8BpmLCJYDUiHY08CoNEKSAzjV4uEyoepxtfle8ajzrsZ4
snIpLLfjtjDlX9Sdi5NiPFVjsI74b9RZRCoL2sEjK+mzH3kra7bHwZTUvgZczqx0sRkvKsu2ISic
3siCT5yx9Eg3XAORI1kdjAanOO2A9jm7/kqY75NpeoSekcAEK54jabPzkX1AlEBWvg1f7J3IC7rN
8hHyhnLQxj/hIA/UtWBPNUUgyXv4rVrbDaf5WkYVV0VXRrs8RM1Ua64MaSih7zFyU3thhxjbdCn5
XdDb0Oel6WDsFnGRnFVpZG3WI8eD383RZuflIdLyHfAjUaQBHqTCkKUFHRwaWX/iaZwUutS40UvC
YQKXJIUhJ6ZgT+mQduvvL7mHm2/Kqm4af3WBoob6Pl6vf64iil/pNwqGedC7bFHcSzrIFPHnHCWo
YmeONB9PoyBiiNhlp8Roz23wS0VVST9U/qj6FizkkqDxYmQdDX86YlGS0T0pVhg/IOCg4R/JVl7C
MrnGhsKMV2+KOgek5bVb62eIP9Dr2D3bY0SFDqlKM1AXBcdGf7qdf9Q3TGVtSMgOfIRh9PWzVHuL
bQmj3uS/KItwPud0sD7dsXU3Lv5fRGSYrZP/Ox15DbrhWOEIVGX1rtVXgDGqmpi1QtGGof8V5CbS
EpUM1aMxiRQJi1NirPP+35Q+O0oTM8mDYM+u8vL1BqJURxk+Lhs6MXWYCRrwH+70w+nM5SQb24LL
qXTexpXKXhWZK0tG0M+ONk3OrQJ50/GKhBmPyOa1i568XWfOk4m9zpODJCJKLtpvczGB1IKz1/rW
Q0JHyhft3XrgpWwvcAYJ3jWA556DZnrVnZxgjnMwPlzIURluoGlz5SN5rNxosH0ZdGdN00m9oiEC
ueVXq/rBP/ivr7Mrz6qywXvHSlu08jKutDt4MS5dguGp1kdpG1GJx3eGZul1MFATMQ1PlpUGJ/t6
1DoQWlSNP5wgDH0R9ahDqIiAF/ghfG5AXyVHBRC+PxHpduId+eBHruPxH52W00S7iDyDWTDYWSFk
+7DdKWRxY5VZiY6qZNJHuK9kbWfc1ApY+884cyhZwBoZ39pD8m5RJyJ1lo3/3LhwtEsrTM7ZS0p8
RA9hwTntb2gWMuWBOxs1Gu93aI4f2GDdWvyj5HfXr7I5tpYTCxC0oPrF1WfEkmOp3Ve26cHXI83j
0i7V2kzmSLDbt7v+XNlJlAepVukZ0vAvDbSjJJYm2SxReXTB8p0K/Ab/Ve5apWOQEWm0Tgdf2Jny
6HVWkUI6prPJnbZJ01+tIjmMMswRaRACp7s1j5nVqR2CO4kfcPlZ0y7NfJYnKvJ/dK2KeLjLpghP
WMJzGP3m+vlNA1Acj+DY9mNF65mEA7rNE4pnshfj7cbQc/Ji4mRLd1FhJu0I5HJq5EBExowZ/MEP
9dlMYLhibhdAqigPsco4T+k3L+pXp8ReKobF+c8JVQnXV6mMKYA2A5oR20pRGzXcSpR/gmfg26Ri
Ehgu3GhKLL1lllHMYQ5aXPMctU1A5ZN564bNEW29oYIkhazAbmFM3TjWffeWgOU4x+J3AShstYDL
gcaqa2ihjB2FQSuz8mZYFKAuH0m6dTLjTSBngAVBwXBo3+0PvQfkF35Zw56zJJVypYocY6F6Ne4f
0Nsh3OETUZkK1vAFg36ub/8lAcHnrrTGZt0v79x0D4fQVaQGMXQxRAjAe7i8gMNEl+Clc3HkpeD1
OsBQelppD3zY5Z+H1wzG3QUiNqAHYLRx/oWsTTFx8Ffv4eYsIfKp9mQ5jrkHlAbHevKKLvRWmHu1
QrgCj2htSmAVB+zaSE3hIyud7RhCgCbPFKJBt5OcNOCEaT+qZR+7TcfCtmAP0cwyC4cCt/C3rcqn
mHxoSdqg0VyqCgSfVFZqlSB2T93VHE3xP2APHlyGcF0gSIcSDEciY4cRAfrw9cVHJTHPpCy4D2El
V7aJtijLfEycCMsEeLHLbki5sMgWMK9xPpVOxR/O7OqCl5WBmJQ+BhGyhWd1UfUluQ5ryCL0ymq0
XHc6CpWgdRpHSCFi9ykVOdDYAdwNSMd1Uou/AytwP9FcKlw8mr+h4w/8BB67sfsBg0x7Gk6akUPW
+0JCOK7I4ToepaCf/ilERGJyEu5w6+4M+qYXAE2oaFdlb0IdR/ldm/TBXekInC5+yZiEMJzGCDAU
FFGqWLbLYQlsljCHaFhcCYjiUN4zTbIM9NGTZR1mw3t4OEFmJ8bLA1Qkja5eI+1Z5pq+rOjXnvdk
MUbWEVb2mfmxrm2PPYrL5eM9XAIKPRPOe5o5ViToZDnu4n2DDW02CsVO/bgJCIaVXlYwk7DosG7M
g9CFrIJkglYsfqq+CTSEQpWuoqYX0Y5uoAx42adzvqP+4pBBvThkT2axTDpiD4SIHi8aYSgiPwg7
AjquVdRNF2RLehyLpI76AUmcKxftZDik1DzpqeMRVcK1O0DFqtPBmEicfbMlW78b8oPPUMS4hQB9
78QkGnCUdNz3SrdYl+pV8sneMWiSxcRlbxysYkEmM0ZWvxWKbs6ZO8b3MKJPZQFNiqI3nEsGfXKo
1awJRDtk8FAUD51zzb/XHfi7VyhTZyoxxiU7v5LA962Zc8AnRLyHoikM4EIdxcM03jCv6dAQMs17
YzSPzqqCD9x8UIyOdqNPY0Q0X/bUgo84dBl/gkVa+nwDYv+aaLF3niI4210suC0sY161vwpYtqzm
glAk3VBPfoH8GWNZknmoWwsxzbxPzoMihPco3/nk3xTDCxdmKisxYXNMdDSqg04/9Bl/dUz4fBwK
eqbOei4CG64FNLyzwRIH6o3u4K/H3XW/uLRV9eOEUnXEzQAG2JpkGhubM7kncEBhDfouqD5PoJz6
cD2S8aL6Ph9E1zveAQyzWwmVtHUT0NeHdn+UZAQM4syFnK+yx85OWM8nCJtTJRbU+F3v/Ic3rval
LZnoOO995xnqD3HKXRCUw6EKl4MVHU5E40aaVmNZM7IbU02ID8GD1Jw4oW+T4fs/oArN0x0PA6ge
FLhNVELA8Vd/mJ8yuzddG5272h9lsNF7iX4OCO+5CYtR8NAPrnkP6Qm+djn7b53YlH6GT1hSioGV
WxWX9qf7THiLrGcs8nvGbr9b4Rz/mmuOUbnMlh3BVam6dhwiwaAccQtQQUPBGpEFf3u7IWZ2k86/
UR40XiV4gbIFazHZbNd5AwMbx5TCGxxoMfK+eRETe+sZwqrgm1k6Ra7Zm5KUZsNfI3Z5CyZgS3uv
CIFF6aPFY6Nvvg2wkWY0/d2dfjt+Dl9ZTDtlu4aLBrywBbYXJmGbgxPLENWpdmr9v5AVviMPOs8z
sQzYJto+LkH0z4ul9mltyG019BgvosySSJsABVnUrsESp6sEI1XrQQpPiv7ymFRP71UJIGhbocGE
WryWy6yllVZqh7eAIXfcOaXaY22qkSJyuuGd0glZEeJc9YSnCeSKjdCOLnKP3vNUVELRNQFo5E3W
9hog5j5bme9Qa+KS3/Ro9NSS1ZmIasBdggFpvDj3kf3zIIYhEvUEIY8ljaxl4H1E4bLnx1RVBbMX
jrVc0FY3xH3gC7Zz+YFqTo3GuOyF518heZXVmkDPlSz6FoeA2oe1WQ6/SpvZPhf5wSJ5fJnvaRAT
Hc6SpyHQDpz65RO8DohfY8K47mVeTWRwXvG/PBEK9fVvuGAf5iqBiEcnQnvQgJ/2dsHbi+AiSjdh
oEwTVMhBZSJprWFAQ5+CLHuuNv5trQAJ5sKgdb9ww/sn29upWcsJSD9p6MFeNS2htR0ahVsyX1ia
aG8+vrjleRXePWN3wKKRNZNJpc6532H2w+0O2YPJ28z/zbZ8I+HilZXWPnONhis9BMLIuC01kOBS
EEtKDc+qFzwW5k8fQNJkrAsOlVsfMNr2xwsv4hCRai4kBtZIRd0E8+S5evw4vmnJTLmQW2sm/PS9
CazorPh6oYMq4eYfxypnhl14/d+18CUHlbQJOkK8ZMxlg2An+zaZBHZpOL8W5LxJ8CIx0IYvO5OK
jhFtdhIo8TAuDi3euz+m1bTuvHoUkuvUX0yqWNwkBZFgfuQUZQf91j36Sae6VANrpFThYTpey2w0
sjXGrZQBiSeiuWGmvtKnmpgs9CW7f3nKGqzzx98+LF/FYa2u0WSfGHXgnu+WQVNzSNAwOn47pPJA
OtmwJb8jYVZ9hHkesJ+h+3XEe5zvIv9uO2OFbl650p0vzwPftgyKAGwssBweh49JcWLMCE/H9clP
alS0RuLLRfVAGF3doytF45Z+TFNMw8wDe7ze6zMFWWjQxkN0ieCG7vgrSypu+S/6ma9Omf+AVzKI
JQqsxTkm1MYy5B2+9qRaJGSxYegULFYHGf+lHp/NXb4k0cn4bX7S3jYEZBHSlWcbApWOW1HX1w02
RHISbbh4zOQMfa7wqT7G2N7gidtP9YV0J6QY+t+yxlxff+rMkIrvj+iGYrIx14ACPcqca2IoxCSe
c0dgfj8Sl/k4kIJP8xR4H/iMbx6dx4VXTC7AU3TBhl1wNS2ic+A2ZpS7P/jPsCAhBj2tJYFirLPW
68zvXkaOK2RYYvBWIznwZhC2KYicr+qcbqYUYFQCN27ndq+1OaMCLK1vIThuOs3MrWSjvYghM4ff
+bGfM18CHz18MGUcQWgO2Vo0goRyY0gU8bNLjing5SBIYrlQvrr3bvJtXux2H2HnUy00xyv2L6Ad
CmRfOmxc2w3pZppnUTZrPHwFNNYkLGSUUwtOi/v+napZD5GPZJFaOb4Lk3/LeeYlkf8XmkXju4cY
YnO7rMPP8lfOv6xA7ZtFLHcbADvUzkPxFvYyR0x/dNlernfXc00kpZ+Fq94UFP1nctNm2jK6pLLO
hX7vOrIs05BwpvjGiwVjf0/PFCQ5y4vz7Nomno3BHRL3UCpYoXU/7axaVxAj9b67iSwmIAqDE8Kd
xvL5dnLkdzds9NxJ+2rXQRsGCphL1qFZyzuB6ghTxtMVSbO0OkkKa8rTiya7wBSMN2aDoWmOQPlV
3PhNG8nqZKgvJT7/nTtZxTTmmBEv3ZLbHKQVOP3JTVoTOBlgtP6hWnwDNt4L+8j40gPhdBanCW/c
HzsBKXvQcqpw5i1ZOIdmhwsT2TZvdFTtUBEnnrSdZ+/mpnMKW7NB5XEZKIGvBbyVMzI2TnB/6r6E
coXbsGColNBM7qDrrft1K4sam5XJcNICNdWpFSdKZThiLPGaF/xA/UEpQDwm5bY+taoZ5N8/hcZC
szFZB1CgxqnvBBMk1FFlx43+b2cexSZ+EF/K5Jb7Hq/NzCnhoHJHtKSusFlhCVc0TZq+vdybZpga
VgZ0edDVYHlkBNL2wz45D+1o6gFdBzgauok0Y+gcINNOwX9Za6oCo2nuKZCMwJTH8YdXjoUg+z8d
wPg315lJR/efMXc/tAWVZX1GFZNJiKE6yNfqaIfZaD/RAng7g0Peh6zV01d9+zeNKv/eiwjcRbW0
7/zSxJe0x101tyCf31E6vMqcgw7/TKLIxUfJw9fa58JJmKbs30bYoYTCQlPLUVPCNqC1UbR8ypeG
FRie+j9e8ntoJVqU8K240zG7fwG5SeNA7Tce9y4sdh07PB5+JlBUeqOZwinS8WmNZOk4lD8GG6mf
CNed+s/ehsxwJ3XcJgURu0efJgEU1IQ/FMC03g3j9KQIHBgHXpRkRb4WOWFqhlkoQaTw/mtcZL6J
8V9IREJhAqYZkgcZNe/+wdiYe6bRB8q5/Zx4cxJBAGxjSxnaYmgqbWbyE+KgOZZTHnc8y9AjcXrD
eBhPkIG4HcTow2nXpMwl1EsfBQ5WZ1DJ7pIsyZngK+cmudFz4oSDCv02EDj3m22SB9JXBSOHu/eO
YBiFSXfjzjUHfQinOrJ7Mgmoqznd9HcQU0xB2OcXJH5pLOgXuTH3qK5yh0pntiGH6borKPzuEXCa
vMa6zP9+bO8SgvaSeYNXiaqt54EZ8/zL7uxHrAuQWeRjsLT4b0MhohODzUpwPs5VPbU2+HaV7hxd
JZuLwxNwyYf7fBRqmh4PoU+5Y/FGUq1RyA8+m44GgLHaUFj5+60PswkRBEZA/ogvPM4Ly3RTyKhI
Ml6ZZ2wXx6cZGyE2ssrEjPOxIzQHCdDGLjWeCrgFoeS3hcYMmfgU4fypXtVXhq+v6E5KiliNQwMJ
nU9qq2z2CvpBhfYWGNlXiH8ERjxtJ6CnDqgKcb1ex4HBEJqSqSxdEEKisfFzHVwePIVrao6suVGy
b1B2l90pNzAT1MrP8xoANAiRAt/TR+l5v/SFRJ2ilPt18yENOOzhFNWcPZbi3301nDYdA2OnViwx
CQAzLIlTkemvAOrNoLJ1Ce8B8rHuzTMIxa8wSPAY8W9OAymxyeiQ51veS5MHaa5dXuUwB5Gm/eQA
ntffVjSF7aRhJsUWJ0gaTYMmV0IlY62OuE4x/jT/T4fLl0x/+neDGZSKbQlSw93IJp0x6dBfgcS5
1GjEkhgSWtcj0WagfTzJHCCx2bWQHQ18z/VS9ZXs2jXnvXkXn2tzeczuUBj4LKemcw2CGRIUwQZx
t4xxJHYYSe29NXDIGiqOteY2nGPScZryawRoaXReD0ir7Zl1ysCyqwhvPqplLKw4fLnpbjeBUeAx
dg16KXEv9sT/47T+I3uWlRe4pAThecfN8aUafGTt0r9sJsFqjaO9BHNl/hWSn7lQUgNbEju3nL12
IFJekBK1wwWHu8AeC94yVoXecHVZ2S9lMbFsXdICYe7AZiI/k/WlzfPl7Lr3k2eO5ubZmAzC9KoD
k9saiFYOsCLCeycuFECZTAh3w/vMsG4FI/HInD2qg02WI7pfZxT+yaNDgm6wsuNKs6uluw33oFp+
da53CiLgD/qY6C/txPUWRh/p01m4AhG/VNTRY7aUMuVshnns3ZcKnvVYFyhAvDSiVKEHe5DMcRLm
9iTiQHMzm7H0hdF09l39psgPJ9oqtWua1PdkmhXTITgc5BRcz5Q3y25zkOydfuWhMdP0sD+kyYPH
CCdqqkA586Y4nmtkMRc9k2VbQj0RzbueLd0niSUV6RzcusCPoSPDNNX/n8dRI7z1ggoq6FF2OpKu
OVngm+E+gFB0aLRnuspmJFu1wAypH399XorYlbOHExyWqP+0m0yMj3MiGFShYVbjtcNu/k7QUaGA
xpCjSuGd38U2wgcg9QaP4TRz5ZO6SCPtaEjUc4lF9LnzNPeyy3dxghzAAdC/S+yNU1SKl0FlbeTI
knI+ADfF3hJIF0R5WTeT7sHhPgo66Sr/RFjz7XJ0SD7vafevi+b1UDoQ8LBlxpdyZAvyXG7TFbMx
Ryv+9IYCjSeyv5GK/ehn3SS4LTqKbbqbNSEtaRsJA7ROhF/YBIJJr/y4QNr2k5A9KJhxTcS/cZ4T
lWeiHlWrmrreMQb4svBFMmldSe1AEIHDxAZynT3Ye2qRndeR0SFsJ1IbRs3KxLTqN3J+owLBpzoo
iwOZu+AoPohtYf27BX1bukIlkhAPg95qP58MNo5uAr/AlN94xJCT3zzT0TJTlrYFgt/k6rck4ACA
kJTBnBqSS/EjCIX+r0ouxaug8V87NxvsKUGA9v8xxgkaaMoEmYLuNWT4gpGD8ixIHLVTFSwpyT78
lDY0uH8DT3IoHIHribcblvzbcMhEejhIPg2ANv/yoSWlpyQwiXYNMdThNb4/qPxRBBvJGKaLk7RY
OWjNo0a0cSuHKl52oJNM0VrjucFsLUAiKGayxeAt5DWMM9tNFdK5ZemIMMnT3Uw5VJmk9/1UCY79
y9bTS34CxqHH+jtVyEbeoIXO3YB6NaAF6BWpqp6Rx84TDUuVge4dXNdbI2wajMp629mhexhsgYOi
Hezc4RXv6KqNgy3NudOB+OGEAC7JaboFHUOufDYfhkWZe4a6Bseq/8/HqaeU9fz7kURRAOeQEFnI
xqz2fTfyEU2ht9ys5wM7K15gIxumnhy1izYoYJYYOy1yLpo5j5koWWuqt+4nwucTnbgPEx0EWB3L
dg+d1B2stj1xU77Orpcv3yoO8mVQc/L0PS8jt5bCn23gN75J5vrl5DjTqQ7aKim6zHdEZfTUOGLl
UJGzQWY02lq1D6XKi15NMp2MAur6ebmp6Qiyx9GrBhfYtjPxgP8wJ19S4zKluji1xcUS7Iwuo2vM
oX023wqVHTTWAzmGP01s5TljpKDAntvA0nI6MHJbqqfxpqdhL/lmESXPVvkej8MH+DprBaaWD7ut
3UmStgwYg86cQKEKYRIcU8lrrwQTyd3ayUaBFc4EdTN385gELoive9Jnv2Jsu9s+ifJ17zJ9T+Hk
pfR2BwaKOlhTFl1UF1eofYynBYGvWzrE6H7S2pnyS0EEIuOVMzTzLJD/PI0p4KQFWAbUpNxMDkdT
ej4/Xk5O0japWZZjgF2EZLhE+qHLEfVB2MD2S6+yKZZxqvCEor+xxwynjDlv/eLDTYtlvzCJ/eu6
e0NuZGa6sWz0t2JwApsHmU7rwg+EHbAgqTYVJwDuZ37Y4PBoOTEVl3BKfWYF7yhaxcwIkVjNgzDU
TuGJmojqfDpOm0jpl5XQo2gV0lqNUvcuPiwdYJApDTzCR6ZZRbDWGjESH4h+CmuyBcUeG911u71T
s1vKe0RkRd1r1NM72FqC8bhmeqqrqbhdYG3iZm//12/T5t6Abg86B6UtN+J3pUCJZKbeqlniVWus
ULpDavcnCZKsyKtcWpBhBtk1lPcH/pMHGgt/PDzHpdYzz4IVxonwRXwZzhPLKCHRZGvY/M9H6r9N
xllaf0/hGJIuKDP2Ul95U2esg4E23Z3gUDyzD09uJQmg4VcdzBtugGAKttYOQcrVR4nv42asEgue
IPIFN1dQJM8fHkzlAxZ+wklL5XlTqtZ9OwOOXZH2WOEtQtzG/HcWKekGdFjEnx3WtJ7cHyv59w5m
r3J+TT6l7SJ+1Eg9upJiICxaYsLQgtDlApQLoq5j4Wy/cDE/+V4RxTAIjz+8XcsDjEd/qJJYsKsi
AAyIOi6/c6i+7phcq3Q8GjIO8T7FXg4fzYUPnHMje1bpGLV19d79NMfo89TY1c7H7jPuK4Ev9P03
iuGhRWM8wxzbzWjomvQaHz2hgFA/MjNe/q3xi9+Qefx54UspAmYk0AR9PXoEO1Ge3tbeQ+2JleZY
cgXOGjO/SVdXRkgc/KQv1BiThuDehWUIOOQDH1YR6DUkUwcjVdt22cHN687DBko+nywdllldihZA
zFMW+sehVTFJ5PoI8545uqqwfEFqVfx2Wl48Qvr/ge781N/c8OG6zbb9sB4QteAEPV4aEW87klkF
RDn7xEidIy4mX92bPtWD61UKsZv7hcJasnT+E0+P427yVJ9WGQhur5mFb9Sg3c+0hlRlkf7A4j+V
0OtSE/r+4V5IaN05N5I+cN9NRCzD3lWCCp+ZI696hSkdb6vXUAm0DN2ohqOdDEaeEzt4wVqKxiQD
TL39j0XYdYkrEOUbQKghNfplRuIBg81yQA/QA41Y1g5BWGMx3i3kfRbBF0ASCpBAIJkKHj11noCQ
A1oOgZLZu6NXe+kt/N+Dj9su6QXnDqDfWirjI++iC3N5z6ocDbTXvnCG9qRCYOnXesxR34DD+xY2
WuKO5lzA1aUa0sys/E3BFkrw/k05yXb9AlICLkdzyWguudPoA066m7aOOrcFVu2IWZw9FCW6ZZaS
NSY8DwxsBVBTGd6MoHA7um6MUn5V9KUISt/XfZzgte158+jkK73pmKilSPjPzLmHFoGIkiSrIDlb
deM1Vt2WX/LZid0GfgIDglMo8sFsqBAUMp44qIsNz945Re/unVdT6eq5SjQMClAMFp9fZ0tQG2bX
feUlmwrFhZBiwU0DiCn6JWFfC0F6CrnEuGp+FuQ6m0KCvyj5ya/TdU7BaoE2ytK1iV6m1I4g40H4
A9OWXVdjKaAcyk6yPHYhqIwxkoHNWs7YdSco6RNjrBPA9vEF8r/BoV0PhLKml6CiiK2/Otru1Ccf
0G7w68oJgmC85GsaTqtMwDfJEFLPMYYk+MEVdvIcv7ZLdfgA3WZt+XojIXp5nsnlHuLIKTe7xcf3
WPK6QHG3jGdf6dJDMKfVsri3J9QUfuicQ00JAZM+tBW00JfqTv4DSWfoMIDm+ePa62k++ngRoFRU
YybTEIVd/1QdA1Ss9ghfyG9SkMgaDptKeDmPv2DkKX+2R85IWaTXiSd5q563VRN2CuGe7kZiCmS2
00YDqFh/jhHR15yeWER73Its7HwCzh4dKy3ElhothQdEPF2VzbLgfQwP4/Inpk0mRZnAv9+fV2E6
zNj191o/2Lpsb54UepRL5ORyj6dWYGd8Iz4PWOCEnJ6AaKD9T0NLjEBnV/8v4X+lOPviPN4gUwGv
k62nGQhNaxgoEKAbzqq2S4uexpNtw71ckFqPbZ8zICw9IkDMHK7j5fg5oTLW8uOF38iZ00LlFjqm
Efnsp1dq3tb3m17v334la2BuUDfDeS8pxEwfm0vaenY69pB2DmcOMinOPcTVb6pKOewYrTMDI4Q9
e1n2VGTlHh0Z6OeDgNqq2iKnTgMx4UM0jm9ecp7UhPeM1Jnhwi1mU80TN7JpLOUATw6YXO47Vil0
8XWyK5ir3D5O0XKke3oeGh1Gybe6IxLUrExBBhZCfUTfR2tMebICPzNqfZ+2pEpJDM82VrtTkyw1
D+xbHdxnpU3tn8NXXxo+L0gKJtwa0t5veLIF3lrVyNhfyR1RTen2pvRjdgmu5E888Nuzu8w3u46f
qbAslQnIjsAbChmfzBx7E4o82EO0o5iHqgjmxfuAKYbcAN5ovlpbfNQ93gxg+cqZLVnOsoOTZh3G
7lUGa+eoQNtor4hqywcpF2o2lKzfgYv4ZPqdlGBDKDi3TpaLMQSo87JSX9hucW5tSmSbGAHu+hen
TXDUjWjIp1oJEWOEAmrJCH9IbkZiAd0d7BOfjACvdTwrwnySOQYGHpfmyNNOMbid3nDcYMtb0/Og
5LLlwDQQxl1jQIrW0mX0NX/7uUkvPyi04zvni3ebRGejpSonNtHorXvavZXvu8j70OzeTi7GzPVn
CRR3aLXtePwWMMWIGwT5dzsCIspssSJaIQfKb8rb60m9VZeLwoaK7HgwDHyAC0Nn8JZjBznQ0WJt
A9p7vpVUHZsZ6z9rio+uCOIi0GA08GWbswIxkuWQqBJwPbzCgbGWNBIFT5MqdWAW8RYZ23TefpmF
aHmj+il4TKIf0E+z7aXfINebUuVAdmvG4cB08N32K2aBoKZyTNhZpyGv60tl8mBYF4sZsY9pV9kt
kqDyPpvvhucpHO9MBOE4vN5PHFzFuVliV7aEkKK5gHZ5MyLbcx8xfZG8Y3+S4Yupufj+9sMBE/z4
LITYGQaLgtTgDOjbNkb+6YzDQ/acMe99gtV0cO+OaQb/alOhnwYVO+j6dCl9321BF1gsPz96lvxm
YTT98L8WMKcxvccHYW26izxG9bn4fgD7cl6FevcX60ArkQjdDzpp9eBWQUZYLDWxvNhioHeHiBX1
znCzWgttTq8Kdm3Ohxj7Vts84JFcgef3G2rr31yoHmckEcR4ZJrnt8GBMVNTTHhBc6cC1IMxafBb
lftMe9Rhlx6Hr2yS86fREEHoVLTKEiM03emO5OW++qJcU2yCcw6I900xDzUL59HRxgE6H2Bn5Teq
mp0rGzhNg1ZTGyhX2K8YitW3/pREqVZBXkZ+7FC39oh1Na/cPKLFmWj+dIi355BXhjhIH+X7gU6C
nawzAMwQwC7XLK/t8frV0YY+4z9oRRGYYoLlzQvQBA1v9+NRnyEAnhnRMVBPs2B1u46xLxxYSwiz
iP2Ks6ixTe3LG8fkd9yOlpbqMyJjC6YiPezSO3ci40jAeTbGrEBZ7T7yQpWTUBI5oLutVDArvYgY
mgZxqXa1F2NbUPYAW52JxreUoIPIBtBW/SdpNvyIDiXegL9MZ91URulpUD8+X00npjhExBsLxdNC
Obbh8S8Aht+cSHQRmFHVKbVcrjWaOkwdefYe29BNSLf/ijub35d9dYtpG5Pzdxc2wdGXeCVomTek
3Ivy9pEwzY3rbJ4Kn9S6RSnvlhSrVzExP8oiCpom5M5/N+tSLS8cnNQz9JpfQk/L+o8k93/2fpnc
tsoLUGi82LcBHd7TrLWKORX0ofe6l26Gm5BftpgSHODSfDz+MCaP24wU8N5iEqEls5smBS5ZNHRZ
9VpwevkvhfDUwT0IkWG1wx/Opzas1OvwIMkY6t/mBbGGmNx7nUIJQo7sd4VniL9W1aODPRk+FdKO
3Qogrv7Ez2AABZLwSgcH7meyxYwrZxvWP3E97Hcv0Tny+Ut7pDE78mKBlWyZf9WrNr7wtb+3iMl+
nv6QBxTmAIu40KpodmNLPyPTBmQxQ/DCQgCHpgpbwWgPAZZHW6jF/6dKrxa4U+8A7Xd84u9gHPaB
r8SlGEmjRGgV23V8jjKAsPGkrEzrpHMXrTLiWwB5Vly0initW/iEZlkN62WJnqb7OFFhZD7XxCsj
0lJuQOm2slilS0um65FIMyMQb3nTTv5kUHY+yNxo2Xb7k/RK9oOaD3h7vpr+pO79NTG+GCPa+uXt
RrWmFmg1jxNCvGIrA92kEau5CVDELoSz5tjzsBMbVi6464xYe5hHUd8sNn4gVwdd8x/sFZHH4EVd
PvMHzy8fEuWYmKZc5zJbPXuArlXo9spHc+CI6N4LliXX3OFR8a+uQXmLL/wAzfISxSJirXCNHjRv
B+ebB1pzHJM88VNGvWc0n3GE0DcWRH1A2ok11t/DTNkX63Zuk1TLVjQVUDpmX68ij98TU8qN0/Hz
LVeZzU8VnCNwU8o+bPZPeWJMxWKRTFHBx9hvfLBFB5WOioJB+L6XcWP78iuqw9hlH6Y7yDn4VYWY
CRlHcVztnW6LaInfxJgw6MJRLZmy6YSwOyfvhNc+9gX+Hb/MYozSLBOxPqdo2TEy9jtXQzjndxQw
HEA6gm+VKyDnpbltWupeFgKIu4KaZejBaJnCpNs4qDGNYLWLqd6O/Tg0HA0p5srb0Y36mDg94Xdv
w1P5LILBU7+Qw3JDb08wr55oea/Szh3k4dPMeNBmRweS/8i3pJlXeE3uwMql5xxg5xVD96hpfHpY
mLULg681vzO3TIwXKrw74lIFq84ioDZek/l/au0AYyXjXp2lOjAZnCXEZ5/XCosTOgnuCUVKCMy5
wf2GSjov0ZH+tipA0JbBn1SpueDQwnVpneFRL1/Vu9xzZD0E3/UmNppMpgvu/aPm+73qVrkbz0xg
cMZjBUJHiyfl0xELneVgw9Yjuk7iTMzpwA9kTrV+1awiSZya42pKZGNhKSGGzkJDE+rycb0PpZXC
CsKG5Bdy4Z5H9qSdzjGocfzFzuYG8qPfmpqLfyqj8xMLuz/SwXKGc8BFaTCSYEsu9Zs1pfKhlEpL
K4gzF+AxAamtN50WYnsxi9OvNGex0DuZDy2HxwTPGWBz3zDJAiQAhoOT0/t54S3EHjXng1iJyQGg
cYXUem6nIAhk2/CNhrixKBP2vnLuZ3s9cNz7VTQvlFqgEn59joJCNhnG7wYE4ol8tSPYYJghEEeC
UWDsT4RggOLa4pjkXPVm+SlfDWp5pFUqeBoAtyo6qG40yfHAA8wPBQLBbGQ14+NpqZ7oLnUlfV/x
WaX2LkS0BMGj3YcBV2dXgVzptZG4guBubUI+AT042oxUPBK1Twiw4BxriecZE+KeCFb07e+iYdhj
Ps6VXtk6jUNcWyLYX5fKaP0E4Tkuc8QHAxKGWOLAbZX4DyAOrR2VVmpFKOei/uoBheRbkILO5ocQ
BBwjZvEkwi95Q1wr2/jQIWRbaqZLfHVv6hbMRlB2j7g8Ma8WvgoQhoS4hoIoCE2XwV8nbIeBHXXo
OnanWzYCcBDUZQyxsvY+dsTmk6h83RX7yiLliHdxxyTKSQ/RMikep3/2lPv+kzkEorQ2Bwrcihnv
pv2NAKmHKhEqFSID+J5f+f15a/QB8+qouN5gorZxeBKA4+hjKfXXt2WpATm3sCtmB6c8+5jsHsYn
0rWOer6HSWJ3aJefFEn0kupvvP3ChIQiydlHkkxyXrDx9qbamfWj3wlnZrE2lixjZslo843jip8E
XWGMLHB535CSvQYP4O4QShwIPX5zCqd01cA8uzYy6uRykCECU3M19TICFlmmynAytnuqU/3GCwpH
cAjqQRFGp0h/XRh+1dhZxEMzr2iWNtDH6/X4FcqR0xHh10JMDuNdvF/zAv4rWcn4Ymcx5J6fiAEH
+a1Eb/Bes8yZ6TwQ5cQN6Z9qqmJMn0SDQgBDowQqTPdm272dWBpNbmHeYbyJ2ffLaTmROz10rpsh
j3TE/Kes6MKwKgDSeupWl2lUVjIT4UQLIlm1Z89IcfdxJ1KVvckE5LXTrn7blsjNMnqaeasRNs7W
eBYP9KlJNtUCHTWLwH7JtOn1Sn0Dd8YtyPr8WQfd0rTefPYU4SQ4N0DK+qVB5HPLt1ZCSGTEMow1
9TKNR4vXJ7koiuQvzWUPPaZtD/nocYc5+AM+M2emqrfO1FS0l1zjUfeYGn0xeBfr2BKbrGKX9Ud2
1IYhIty6zcYfGrh4Si2jIIaAY6jRWdFHFPQvV+tmqL6OKk5Kr5NTaj+N0zqdlzX/fmRsFbVQ0zxM
6qcO8ncOR+Rl2wFD77iGVn0jxg+uLANVctgIecRITE+l15SK7J69yVJoFjGTajbNc7mB0USLvOzH
7vfFpEG7XhjTN6fi77gyhxDXY8zTmfjrj+tDPa0TjF2NGaexSNntciUbGjPXq4P0YpdbhuZTT5Ub
dYZNyCAAtxqojUgjbiEAUeuCj+MIsSCacSxQ7JihU+SK7DOiJIG/WDhHJHQ8sh6UyexzgKaZyRnK
Hpt1wnugzGYsESpWHptcfSfIKP1rKy3Nu5yaMawOuylVX/+wykTFigkVQLBsGI+24YQKgWUHEPJU
ZU9RDQOyoN9BlCAVW/DfZoWyoC5QIA+iY5KJdgnI+/Z/LoLdJkJlkqYheT3lkl02HUFUxz/h7FRK
GYK00Xks5lCU61yTgr0rw0JuHDKBT4fQ8+r1OoO7zHb358WCmmrDiZC5MLduYYj3GR3RpbnxcVrB
Cfc8N1CUKdKEWtt/SXmx077dAMoshP6kdGq89gfXg9HHMWUsD756pER+YF3gXfvk/79RoAf26gqB
ogTLyau79F6Xpgl5Ig1lOAm6zAidnSNCYcyWv3iBFbV/415zi7W6XKPKb3xQksCCit7SFRyB1I8T
S7BpJOHOb9F/iaMGbqHoc56rrUEMJl/D/4jPYl4GgS8nD9WX3hzGIMv0ZKKcrdAS+C+ynEw03WBW
5+ZTbTFHmoGgWleTEvQY1f3C9JBeh2caOXh49TPqZjXlorEfPTGoIe26LpXPlNEPB1n80Y1hHWne
Jvdfg9lpP35y3kyCJHvZ7yKL0WbX4kkz/f12WQp1YsJ3mCX5n2tW6UUTt9hEnmJ4oUDHxD5nl9xy
b0BNLDNR0USaEBJkVIA+icOaADGlH6dLqXsHCD2TRt2b8nLNKqu1k1H8YOqIHwGBCHO+WoUg9eYA
LU37y5rsJ3HOXOcRKStveOB0tomieLDEkAsp1bZYbIAgSFmb/in5yogaeynSG+qBifq6+jRwrDWt
9U8y3PMyPE3LIBwYSWUOkXQL6OfQKF7GKb795hgQSGSPTiNoFjQU1VzeDbPu8kkqPV1qCZg+W7gN
2ddOi41Tsx43GN5nTdth700z59pBNamX1i9dzSuuW6uDU2YdVWU4y6raDbm063kvyf4V6USmQUwf
hwiMxOj0/pKjg97f81pNDHxmzv6VHy00/NDRtSopGky07BhcisaaSM3JmW7kX70exwxZQEB6GZ1p
tNideutSizx24xegaOft1xg0IcakaF4NV2NAFIP7bLbg14arIrf0JXw/HXS2ElyqJsrCKVjj3Dwo
TWLcls9bMuzjTVJdV+PDyTid6ccbI4nyPEd4OQ5AV+WGaUQAeH20IQ8hVF+QWqyUgzArkj0WT5hA
Ivv9xwudnFLZKF/DIrvzv/b3tDOcRJgPphEAsslZICJ4za9rXQPsRITkGOnyzdl59oaLce5EgZdx
UtUSZHEw/H7VfZfjq0fhyz6BwKaugjUZo0vbzIsaS6XDyEpU6DOJC7iJyM9U/DDBaioChN4r6HjJ
T3XGvqoW69MKp7Pz3bwtutRRdNB61WJzIHtMPExb97mKsNRJ4m2yeECHMZ31uB7nDKt7SnNSm/hI
9vdL6oeoIP2R107jWjdeuY830cX5gzMIpoutr7wn02yyCDePdPVjZHkPGAwcUOvNdZcuuLRkaIpK
hS8k1LXaOlnRjQwF4Brd5w7ia1+baA4TJQJ88yWwovDWbsn+2VO1q11RVaMfR0umA2oYe8gxN7uw
Kt/rCVPCMwNFgR7HR7b5cuGVPi5jNSI0hvBalIFlEnbDdJQfVOaLBO1PSAVdBSWH4KyyEu9ka/5S
2eEU7LVKAwXB67QtOw5CxWFatMX3lr7IjX/WcG2X6rWSkp3mc/vmdy9XBurgvcmL5vR/Rh453vZL
vY6/INmFXY9uQmK+Q8esJm3nUS9Yqkr0qKxGRQkhg6huAzmrGyEJ+NmBkIqev4EDFuoAKdvXv2iT
ZGp/ZLf8/HJLSHN4SQLn6/s5jJedq2mWFnmhZSktK5Sq5tIw9QnYao8WF3zW5ygk87RMYxfU3vV2
SrUqPj6uUb8JtSK4xktmCNy3P2Y1uQYrsZBGenWkkxh0Abb1IdYUu/K53TEplOdOqLZcBNLQIrtw
ip/rCqORtjxzA7Q5vcRk0tfsAVHWqNvp9SbZ6iGP4r7pWV6LAT9k105l2zNX5eb2u8k3sJpcBfZk
tAjCYk8AjYOP0ggXTyefz8W9XADAnHREvffi1KgPXoomz9k98Oc9PZ9Czw63RcedIf0II1P54XjD
2VawxjblVa+C22ONTDez4ytPolJU0Igis2WTnX9bR7O0mZvNu4PIH5RMJeC1ACxl2jirT0HolWkB
yJJChBgbpzV0Z/NB97MG0M9hbvp/sljbDrBsrRYe7x5TM8Lofao09la6GEQ0+m9/iL1HMyeT497T
tSsGSR4DzcQ2znV/or+K17geq2KZZmg8F06GQbfnlKTqjLCewjAhWseq1XwyrCBu2MRlQN8kxJol
vp+XUlpsOzT4Q8FdTFgLO9uUmwEgiaLl8w0jWEhTONpP8XBgA22NiGAXd1I2Dr9Wznayb7XmV5S4
JCwLsKb59bSxgrxm31rAZ78Cezmq85gXpJCNL/wlIu/G/MIsahGcHKZLiV6+VbPtHUQBB5KfACuj
iuL+4vyLWEbB5YL5j8iLRIlhIf1zlNac1UGEh7mtff7SVe09ErfUcE1dSPTi3s4G2TFkhaOcWdt3
n1uywJnEOShp/6xCIftnk9QtXyBvI5q0BzhHEsRMh0YjNzd4dS+6JCpN9MYGit+i0io23z8V10rf
WWH42bJocrPU0PoQ01m+lY+bAK8TwoJUjHG22ZI+aOoMwYHD7HqEXHtE1BZt8EdvMWRilzBjfVBL
OpMjztH0CPBS9lKcd042GIwCtrYSPyvcpwRN4XiC0tB5qEnt3rf8OEGCkDrus6GpT2eKT6sZt2eI
bn43OZRePyyAR2eOMQSmh6O1keumWOUrks+DxOqe+2603TYn+eLrhw+zk3/GUR80TwG5IqVXGdtp
bY/wN0L/pzESa5nHR3gtMRqORNVfZCPxHPCbphmF07XjTEVIdwBTKELpTsjqfAtToA4cwjzLzBwf
Z0FNNKi2g+IRd8fTA5PIH2cs8KGvbrzVNwIYVtN6Hk0JcCIujeaJ3BSdx1/u9x5y10hYvboGbIHk
UhCG/Fs6nJr7REKZs0P4zWQfmLT50Mo/OzvHPYOx7/1B7WoBGMEZg32vKcYqxTs7xZQIln5NltZV
1A8rrVIYS8TgZzt3aIzLyRpzip2wFR4WwxIdVRI+r9OJA6URiXgL0fdy5VsXmPIIwFeQx9j/7dHn
to2x7SiedaVRhXNtTvK+rokDkzr1NJF/NTc96hLhjtyUS5jpxWJ71fnFcWCPY/o7/kOGTPGVyAA4
q5PefNiYKKee12cfbZPVSRDXkHXLCBgm8SthuHFrT/Oog/h6Dw4ZwBJwYNetYfzHJxLQ/K1aq3uz
I271jMkgl/xS6DjCNwv4PKvaAe11YSlxF7hCEqavzem+2n01/J1aormaqmlhXWXTarsHeGkMNrJN
McRc1h+tna2kyMEtZ4gQeTwMr/5RsWjLJti2necm4DNT7e+8sAoUcnef0KCRNPoOGKH2y567QUwc
cjJk9xWW+NF1TjsUTTfX91pacfN9y7fmUPP46qkX4GoXPMA0mTu053lDfzRT3CCnOHG5IXbWsYf7
OAKlbDdMKe0DxIPunhRnkJNPjHHa+QbYrUSi/Zaq656LlwCrhbBf8Ely9aBpRxZ0t9o3btKRXsa5
ssQr/cJ3EUg/mT1ndRlhTykMn1ycOxDGQL45AfXoiLtLEi89cWHzxlXh0leALkkvUJyne/d/Xu1j
Qostz7UGKscguublRUbIsG2sd6zX9JV+X8+1KExYRz9Q+O66v+hFoTQYbeVkR/Qa9li3Y1q8u8O/
0nM+JmKeZ9uji1bQOY2jQFGT48t4hL/kJgk5YGdXoRQ7L5tuAsUpPjTsyZUWZ/HqutHJT3JnFj3b
oAeHkkVHh7zR8NgaJHgDR/BQ7iDtOjLpWi+gLQqWmamQmmosst16UcKBZTTJZYG6b5iUpLh2rr47
ZgEZ413VOINsTgrBoacc6apV84sBUt9OjQbRh58ARLqIvO/258qc59fJPx71/CvsWlDFIhNUcqhE
VbyGIo08tKCiTsi34LHm8cjmf6cASFWkOJAibVtnuf2nkR1nClb/rL1JfAjPvPy9fK57fUEnHjzv
Fbo8WwSBqBBxokwM/pfjmUUxhEsq1iRLbjZrOH+UNzBa9bMb/A5FFHxhTFsUvopRlu3DsA6T4p37
CTmbzBNSOYwF8sSJkO3rKsFZfxldXLtJqrgXWd3h4/k0Lh+EFTPBGsoOtvC3zx5Em84e/pxMjTvv
EvRFZkmhDJw17d+ABKDZlPHblylzbh/7VvPceeHKQyqGl7S5p3jjrwdAQSL2Xu/o8n0bEf9ZQjG6
a22mvHdNMl3ZJwwI3UnyYHeIBH0gk+w87tEsUlni9Lr6QH/OrScagSuHyn7yWPzoGNnRVDhwFVeN
BsGYKT6NRQsgoCOnkCASETHSkxQa+1p926jsy54s4dHgemmmzJzqLIG1J9rQjC97XoinvwkcVy5J
khheh8ATaorWkgqoFMkjfZ7bVa/xyCkmNwtq8OXbYZHeAenr0+WaUEi5dHLZnkWuaamRqfdQuD9o
zN1PbAZqTDFuibCsCEbhbqIO8k7bpppx0sucoF7Wiqewiq4HZN8Ca1LnfLp7jQ2RoudpzZSX7bw3
qWqPWTyH/luP0pC41k/LElbZaGqEAWVX7JOIO1FOn4z6OdKYx8f2b+zqRm9BbQbGG5MSlfwQfOLQ
dJtHeGjPI+a4QQBU0XR+U//j+L1of3NzOnc+Ie9vPYPXIDDxihe6vCqz+dQpISMVG/3xUS7my4h7
LZ8mxKAPNlkvXKIK/LHXlcT5d8Rdusd78FDviHHzFOIPgfDYFenFRpA/T3Xqw8E1CR+WAFs+GY1q
rBv6+HV00OJZ1rXmOqpeHnFB0hTymRSgR4hKsY8GDsyBnXp2r1t1P1hFOI8uwOV7SI4vJni/dGZi
/hslN1TcHQXruBPx992uiFJhTSyqaAhsqBcEnKMI340rcbgSXdup3rWERILGNtLjoz+KvtYzHDW/
vXbRuOcL34BEOK4+qNI3wPOLt+2Nc14gWkay0kJyxk/gss88jxKIHlmsjMEAM0EOnymkxPKg4+bd
YK+M1zlvIm60+WtysQ09iwqLgOxOLv5MuLKu9Kgib5jMkrIp35l4CQk7bjGi70ycbhDgd4dfDuJS
U/qLkkJWGJ8HWKwH4C00PRHXDbHyHKsABMwyiiBeSLECw1ApIijK5IavtW5XeBIMgT93VfNkjGhP
q9YNPMTZhmz1QqWCNcMJgUeMzzAFdniCxPtP/1/HRyKLB4fHd7ik3XXrujEFcKB7eaN28j0taJ0E
ZKio3566faLVgPrKGqDiViyZc5NsLM1Z+pUd0NBMw+4Bp4D1R0AWFuknrHpvlGG34Uc/ZlxxBuIA
+p79jWjJGClFiWQ0LDKW+SvgXy+yfZzSNYADdWIbCiaxOmvyqBRXstqotODpt96kqSk2G6EOPvgh
4fkQziK02G5KoSe3vd8KJklB1QUKC75tfa2b8cUpoxitspwE08RefTUYUzxqLXXx5FT3ZZ+8qOH9
FXv2XbwlJS1lByxfl+xWcvnnMO46Pz01J49XwvYiepaJdy+bld4DMAcsdHuGr3rpr+XgpZXJB75c
VmyXEDAAWIH8uwbwrFx70BL/pv9IQQc8omRqd1NFL2+343Gs0nGiY3/gbOHyS9K2J9JLU9xKge5d
iRxO83mc2VOx5OVUcEZolQMO8+dTWXnuifIzsQ9V41VJLrMLaXGsCgRFCW6PwDRevUnT0xLkSr+z
mEAoxhstoLvPIIfs695bE4FVALJBSf+w4s+F1CszWcAVzd/KFZtLwxa3rF+NkPGwqT8U0kzU/6tS
fk4KFAJlzPhmve0HRY60rZz/P47eaR4si6ccI+IcxkywtbB/iNnFIYZAhOiaP+tV0F36iobH0iR0
ZMpaHWLXrY4yuonkyg+ky87M8GCgjZ5YRxHz66L9OKU9QcWVcle2PnCj8j0nQv6+OoD+boODidQI
KE8OpbOKnHlx27kFQgCa1xE/eOOpxtJmsEkQrcUpOEBNdgg45R4JSxJbfibytMEh89yiyx5TE8Nv
Co9auQIcYLByxgR4yRS33t+i4bqEB57iYtOJlVIeLxpPi766JT5lBo7HFFByJ0iFOLgtRIqqHQ67
HuIg4ffVvThrx+YkubRMgydqf6WTgpW03oyaYM2Y8Ueyy9uShEN7FIU8ToKg3o6YllkI5UYvICs0
9AbNV4fMzW7+lRKlEa664hCBmWsYY4S2rsWJzx7iWv1PUwFTZS3LrkzPsJ37acdl5R4e9CdzBMwG
V8FsKoUA60mWuksiW4d8eFOd0NBXLZS8gesYUqsVSmivHm9TaeYl8pmIfBwNCbGl7bxUrpSdTs0j
fColNr9CnfRnbraMF09gsnUk2cAI/5FgViALy/HDxIuxnfkPcRY0NbWraRWm/9RgMK5Btil5c2ZG
sD245Bk0tz1f+ulOavujY4SqqYGxiLEfUh+BTCaaOqvesAHYfw/qQ8muBt8oEOdV43hYsF2IWN2J
cjq7mxkCzhIzcdh/F6Sk6U6j6R7QZLf1oNyF7XgGQA7VG4s2R09KrBYy5QrsiSGoWc0HaeuwIPM+
nTAXkayWlcn49bgUVkVFhGofhUB23f09lu+TFIPpPBcslquNwx161CbM0AXZFyHi5xb5gpUfj/97
KQOk/NmO91ARxsne+uuxdiINlyjCOszk0viqae3TqcESIqWhDxmWn45DCEjXtDDyvywZs5+VzxNi
2pt/098AQRuFKNcJeVKdI1GjlyTb56NL0uAuk1PP5slDSjzcpGDZLx4YOOwgeXKk0j25nlr+s3T0
6heUvuZjGnI34EFRa3C2Puv5GXmzrAnIcY3cBX7tzXolpYc1b9iqX2hgeccEkZsTyZWGKCHgqpAu
JuUfBObN6QCM2PyJ31mWK66J4nYF0BR2MvK01efgM1/LWU3jbI29RRnGRTY363Z059Yo1JO5FErw
2WgKnOg+6UZwaRashdkIjJm8TCOFzzCZYnAuWHIsL76a9dyF7Vw/vdLVYoQ766Ceye0IN/UfZ1w9
dYWosuADe4BLdLsHO5ocJW++81TBqt+3Mekax/ip6Oqu46On+65SQZHWGe9LOJcPXKNqi3Xkt1GL
jjoEvxGLk/XFcIjexWzZr0Bo7OCEjsEhVn4QBJ92baRMXRJvcEaD/YygjD1eb8SmJmJs+UgVizXo
+1JfsXyAmMEBz82wkebZFG6Z8ghgimWiWaRM16blnUxyQbO2PJljZqS7FlnpQXqtfilZk8bwbe1+
dtEcO57mb2ZKnYBNSxUWQDnOHQVWt1rb/ATfdFg1y35QK4wJgOQ+WJM0eXwOGFlzQY9RVXfLK6Hs
EA4/u66rLgjyEptcx66lTLCg+rpzmryM5IIX1RP3X7YvH08psBCol3MVB5QDR/ou6s76JHXT6kZh
9/0bO/GadopLJ65oyF8lygvZwh1T35ZrQRK5lie29yOtk89ee9sZG8H77j+xtc1/fDZUoWdTAvZL
nI2REhtXdMAaVX1rSP98rTczxNmJAr87LogavKVJ0JaSfX1UNWP1t6yHE3OkCCSHG/EV1aU/h83G
tAGhMvbU/ErBsj4PU0r964DtV9dsGvu+4cCcL0IuX9FjodMtkOR9YRWs2RO8SpSJRHZcG1M1tI6k
euN5Hjyz64Eo/V7Z+6NE8+ieA8r21fCDy18ELOcxvLvDWRURzq3ZjziNd+aT17bDdWBj5oaVzHIh
t61PwDy1ip38CTQ2L01cSoGBl+NogwN1DjiD+dKqBL7ZSF7K4JMU540FyTYSrK7KieuvVVpXyyJz
5kcD7DzUYfPTiy5xTPsacUcfhZRR+siFPr6HCwmkr/uer++YR73OokO1IhPOqMQaUPX17sOsOv4g
IEqtjrfMmv/Fww5qpO9Jq21hGhKt4lHGF1FB6ezOio/SyIKP6rR2dasod3Uw0K+GqY3RdyUaFAX+
HwqATLcmyuikTCdspoBaAFw8cGjsC1JdH8GaiIkdCZ6K5EEaHnJth0Pm/qK0APOzaPKva31hQ6lm
iXMq/BuTAX5rX/9XwmazKAjT6qem5ClHY1AIFag4V+CdGV+tETuBu1Szw30dZcOUkai6Sp5NJ+vN
8VATt+DNk6vDumFQMIJTqt5UP5bEdpweuIGokjEZvED3SxgmdMJZ0OlY+PyQWE6HBIowG4qJNqlF
t8JpxC19gV/C5GBmN5NhYwn+NR0d0Cw2WqwtaNdmNEKGsBm8azd4PnJbdlFPwgWrsQijYN21FBH2
n5OmZdOR4R6ZTqMQSoW6vtKj/IfU065yOJjHk/cI+/+WrKj3pFIMWKwyk0Z1q1OzhkjnyJ4g0N+T
b3SvypaQitcYJpd0+azyreGDU/H6UdiSz1cE005OVy8rpFyAxK0Lj2+5/WU7BIsWf2PLbqdDb40s
knCQ2MHkSNZ/9Gf2yDb0LUfPsCqMXSN3PTjFetxBfTIjl73mVLnds1Ol1GH6bfow9f5x0z+PA2yJ
to9aKJwC/v46G364v3rrgCrpMdnFKfYiHIOfdK9xZ4B7HES3e4xkRQUNdsBj5rcuMGsD31aMvk0k
PrCRFy8gGL+UvxOlF3j2CMko7/HLMpunXkPc86MUHj4+O7oRET9hS5AF2W9sKnWm2jWq4O+2gIK/
LDBE7Eo3aW0u5JKFO3lAhn2HBg/r1OO+E0ofDj3hd7h/oPMq5ehrWWlzmhAh1eWEdyaYE/G3dZ9W
Y3abV9kgScXIhmVHyITsaWKD69IK+ECYUcqDLRvInsaYxSLEqX2ryzcXCxzVJQiplvj/7sTA79nl
m7eOYW9hmD9wy9cQjGxXvt5GPzgwx/oaHzXHGI2E5/G9qeUSdbflujAk/JbEws02/m7eSZbEaJ4m
HYvfsBhuursbsxMmQpEq/4jHqMtKMQ3KJDoaauyKAdBPMGuq53LMJsxIhnLckfmiPBctL/heDqrs
veVoIdxkjUM2yzgzQG0De6CbWP8vR+9F3CkdfnH1n8f1l7mzd6p+81Hfg1ojhn2M7hQG5I9xubqk
+C66EIVYhY/MzudqBdFkzTBXFTeXgjZexgNfWWXbi8Cc+OBM5WZseJSZOuFf9Hy2JqBd+jq0ghmy
a/n7Qhu++pvT/uQ1BwLeFU2APxf3FcNwEtB2s+7bx5k9OeWQaFQz8NynZWHzoFzG/Q2vTaiGWQTY
DXaMI90yfy23JwbopWmDWQPKjtV4E1BEv/VcTN3mroeqfqa+/qHr4Qwm/I6TD13PM8uWes2sHlr8
ng08Aeq3im39aPbp90kqVpgB60x62H9M1i0hiLVTHSv0KhQOSBZJrz5nbyQoTlh4ifq6LqHLqdHr
cVUj5fig5R9tKqv3aXfkYAJa0lcHjW3QEKKJMOPoMoFK7haPDRR12bwvzf1AXPVvTGRZjs32VjnK
3EkBqgmV9XDtG52q5/nNWmOqV7AVUgi67XbBLNoMxqK3zVShsuIccAVmB00QlTCrNbfP2zkLq4WB
SInQ3asoy1paGyRKjooxBCjx6eIrdNzJVAv32aCXBQVnNICYw27Hp5p9qTLYUJMxfyeZFNZUpJUx
bMUqwyb3k3YS+w6Qbe2+qqdNt76KIZwP7QGZxXzY19lnmszMGcuNdpT/TculFL4l1RjwTWrfrLiS
8jUDLGGREpJGSArp1IdhUR/0kIPp9BjeWmOhBT1+DLzdeb4ZlSHKpDoXJoeufywPrRJGvgA6e/PN
fhRR72NcL0UDKtnUJxZ0lETxtQrUmO5iYM9WynOqsFDQszKKrh9lRPUzh3vueO3Je8kdwo9UkQNk
iYMdro+hjfut0yb425sOA4nzoMZuGV5vZFT0POv3Rri0fW9uwfDmWLbWv9XYb9RQ5lrZeexWqDVw
31c6pBJTHdlUy0GPYj1FXNHCKRXVFToKyzTj5gsbzig3YXMhWhjAA2tUyia3jMdUaQhpfVXWNOGj
hsra20kiuosRu22UcEUiV7aUMRIssHST3f5QTpxIrR03YV4EZes5zM94S4hflydNVnwgZaYlenCc
QO0locyZNUl8nNJcwEPgkETs5PIp2lymAMYfTdjINvfVs0HjyqsreNH8Fz0/zFszCMkEnDay1O8w
q5GfHbeYzxNjXcJ7zfTsydEYLjd9Xd0YKZKu/xNJbeKc5L5kZ9SuyTroEyv+Mijk0OBM5uAJgiy+
HevbOBFkevEZxW3uvWvHG2k7dnuj/2EJls9jVLesQo6K5QaBuv3tYfx9/GxBxm80TqbR0mCocKfC
qbhalQf8skzh9tFpNp1vpluBT3GumUaSROZQfH9i3rqZRC9Wa8GEwry7lcIu/5o4cW7Q9MCR81JP
xroqE44sk59spGEsSnWvvUGccx+PkCFgTKhH/PkqRZcwfMEb30dA5n4fufEbTLp8wxC65nOGKNey
qdm7f8wRBWlzVsZry0LHvqD5HbsGDGXc6pjIM5Swd1TkB7EmylBK+ddTbtVe+JuFgbUlXYWswhrA
cSZfPXR096nABn8aELd+i5226hioim2nMA4nGHqod0ehT/OIlSflL43ijtwFg/XSt9nyTndKpNwD
Eim15OTEppIw6Gk22ssLdVXDMY83u7Xxco+GG17MaJMXZJZZsVRA15POBIZSo6De/0xFM1Vi6RTr
pPgJfv6kVIkgOlcTV9G5EFWeemEPcdv++cpJP05bIsmKrb+yBTc/lGQuy3fFu2eCVTIDiGbK+IzO
cVDU3IWJ5pRRUt4cP3rGeIl+5iaM0xoIVeWRV+8W4NA418ekqoel2L0JODM9JbuwakTm2ZIp3U6+
H67+UmeewyVIcsclY6P+myccWJF3m9z7Merp7qAwdgCHfQ5NC997FqXnvEAtGExvQGW99/RaHcRc
h3QsP7Zois84PXadjNN+sADiuoA8wuLqemkQp+wJxuGsbfuhjV32T2utaOM4jbu53gSzJ/x5nici
QPP5pk5XRpBtBQrhzQx6mFT96s4WGHrAap0BqiiTI9tPb1LhRQkVNPrQ09yWBb1feqnbxQSeT4z1
TIRncxTqJOjp3bwecKBszchr6NnkslkXNonEsPHCcrpY/2gqbaRERXNiE9V0I1nDGV9OociBOCQP
BdWFuZWHWv3V5eiHkuUA8z9ZwZAqAz16yZlXNJJO5mPyK+HnG2t01lNX0jUH+PV5uK5KX8B5MN9r
x9VKxyLhC/X4j5s8akCtamYQUNIEKwLkuWbznDvRXSg1VjI/ogYzVMe5SEN70yIChsHv/HHo45Hq
HZU+0XO4/qklFYAK4I6Gr86JtNITdX83zYxr2PEz/zP0BTfV0aPJSxKZWseYsCfZBDVzoqjqjlt/
jOgrgfDgex6EavdHFo/BHlLlbLUtkYVNWplacZovuh83TtB9izlpRwlVzChbMSy3lBHJNDuPac7L
jeSDZFTDBtRwx9DgbhhChNaGIzffyhxKOvsFei4chWhgGfxqjqDSvU2kNHW9RnFwdPVyohWhmDTL
meR+Ol7TXjFlGsQSoAOfZbUiIUZWpclKj4S/agGisSiuUODvRwlX7AIJyXFe8rk21R5AXvpqfnuQ
c6vsK5I0QkF5r3rb1y4asDAkoDT6o0pGXP9P4iFNMDYXQWVZgLrcvJQmRrbHkIa1O0/oHjlJ1H3f
MvGw7SDWrcx8ufAb1CBthfL2GHjV5KaXJln06naMKoku+Rt0VszvnR/q0gY7+WvDPlbdmXZ8NZrk
SvwdZjvEvXLEJChHAcQIO8HSZxUDcRSfUXm7U7O9EUv7bl+gCdBAOgdD5LSc0iXtbcz9RUZ8/naP
fql33ZD/pR6vMdRKyzjQ+Fbg+CbDGDp4agxkVmy1Nk0Gk7NhlIPW/AKb+vzZbeoCq7tXaiJZCDE2
yLMRYkZS1STQfN+Ik+Xfa1Lrim+YoyO6segf318P+SMRQdX5LYcr6+MJpuoBYd6uGfNC12JWBc7t
n5/thr1Zwo69ZUMJNn54DIN7Ytk2oVFwR6f71McpDDsgS27LycvBnHu+LbzLHBn35CytJwAXZ4Ee
en9m9quZ9KNwKkTL4Ms6xPPFHhA2OjEvc+9hU04LEsoRxyfP8Z8W7XeXuvMWdmwQuzUBzFZFFUN5
Dz3hHvb3T7XpowjzXdPZIldQRbdjPE5/oV3TeKILW+AXqpp/M3zC8wGO58fymp5ew2B4k1nMPnKV
jUYKVxr/gFwDTHjlIdKM7KtIDD1xXEJdnyQ3rW8HAHTbv6C98BqtPdTmry1B1W6XQV2RGVmHaSIF
PnZzWZzSjwdDCpSRuwD0fKJq4VhUMx0wiQRg6w0BTS96HFa5LluQo9V2dsUEg6hYKAbFp1lHnB8g
RanWPiWF77feKgdFIzYpegjQ1hT6mYO4PMfxWIJN9Mu6zcQEfBGQh2MdE7uigBZgqX+7I9wZfFDd
r5rJBWJYxkbsEE1At6c3edUNzEHUimnaFPpvIOPCWR1fVmjIvgqaBp1COzmRTgf+Tbj02msRhuXK
OG167/rFEKKXKzEoZ2F8o8mwuHZPlc1RVbDL4sUdVjQz6MiCBhQvjcwc37dK5/lzBpbu7xuzXYsD
t1B2KvOokOwcMJNldiY67ttj4hRDC+zV5p+QbSWuHXbUgQyDEHq2RML9j2JRDyjieEvu09glZohA
N5qFr9QTIuYfAACsUKsG+CX7J6smgSf2+X+E1Ud78fy+aANLUwaNlCWP1SjBRDBRqpm5TO6hHEER
x7Opmm4x4yRFgkBcCpmTB9uUD9LMA/+7GoCSYId+EKYfsPa1/04OBJB+NCknKciKVQlMuwMF5972
ASGDhvL5sLnFpVEbdRqup9x+WEbOjiOvOS1ZwMq876GIxLA5NiYjlvktVcZq/eidbtvixXZHvRQv
Ezox1KBWGZeyhziosPlUGEqplNzShjVXGf5M5A7FKbtID6hrMDn7O4qeXRP5M3P0pC2A/0QbhuJe
ieXCdRivZ4bh08JevI4EpdQ0D9OLhStg0H3+dI1X464OJP3AJy27+gn8t+7XELS52ftFMm1OwQTK
ogrGQkj61VtWjM6wJ8UsUX1UQryRZQDSrUT+jRsZq58NN43fLjjuLWCvsnAb9xNo/pGCjagoECT6
yHVV3oHuCC5V+TfSwXgQEHbwMr99W4fdc+tAHIdCNsRApt54Ee4FfuE69aLAfku3rcjP4hdma/zk
mSZz17542pFY4uL6Mv8qoeV5uWjLsSJaiCaM7Ky+zthCzh59+RyYiTsO2QZsBQYGWCKXGAJVEXQf
bJAzE9IQDlOJwNlvEnUc/gZXrPdyNLTOy7zWpwoFhwPzyr6ZEpCyzbf0sHEom0hK6JEFZoJwdcaa
4vqU1QP/1mnqqPvXIFC9pae6vtAuVQ4CWKZ4sVhzh3JWXW6DOfohrp4L3oPlaGCN6h+tPk+amvHh
jW6v9F68/z7Ew2wO/ExO4/EOXrtHIlkuQQbFF3DO0sHwdYC8euwhKHCScgOH/N9pWm56bTlEdI/Q
D4Q6c0cEceJar+2ECzNnmffmnERrHXlrqrD6p/xPI8PRvGyAE9M8h5oK7mQpEgswP4OhkEZxRWTf
0LomEHupQ43S4MKMYvRBh221F4fB1qDO3fDJETBMwF8sV1zMvFKjOKDpecBvi8+869h67XD6uab7
JKRBnGzxmE6gYhOaol/yZluOtz3HjKcDiUy2dH73CTD5EN8jeQtxYcyrNA4RFFhuv2O3sW+U0uZb
TOzKdEI0G3Ow697CyH/MUfV21PzSS1gDBS5gQq7sbUlE/92QScTVgEwnwWi+XklhtUPwJRzgr2+A
rrByLZ7I7zHcJCnqwU5nD9xYD6uBBRMb9xphRqZygckv90zeL5qA6cZBjsXva0S7kiNtJIS/ISSg
a9UMSbW9CEaF1qKKXvapO23pfCcGFolQAllbBKbJPw7aqjyy4VcPhO+Jn4S2vcVxT6f0BWT16osS
AfkAgVtUgHyJhpGvl0zG2m5e9mzcWON7dWGMyf6sIiQJ8mQ1CgJe8zZPUHNve/lUjevEFAJjGvY8
9OMoY4WfAB4/5jfyVLnOYmiZI1XJrtWU3BD6hQFZgYrVyshKqD44c8p0AYgtMEDsGDSt/YR02Iy/
MMjalKBK8f9uZ8cMakis2DRd/q79iAZqKSG9J6s5bx9EHLUHVcirz2HPmtDsXxW3O3RdlMs/6GVA
hulQ5hh0YL1lf2PuaGxTTOzX89LZKjidjpcdtP9H+b46sKaNI3b0ZoKFQY0WOkfzqEAMM8zzBgcR
7k3oR2uf0+WFFYAbOthY6bxlQyUgoJUjfiWkaViQl0gH00vaFVBR/RJrTUHGUstFBVESvmHXL7IB
HGMTroGSf0HZx71Lt4W3IRt2zkdx5sQBSltB9OfOqYE6c95Gd/1t13fkospkIUS20EqKZyQz+Kgf
j27dwfAQWUMqvE4LvIHWy+5+uWwTGtp1Dq2ehyeZmwCjqK4nkv7WdWgs+hQZVhjKae7HmKGvFy5t
s4Dsxv8q9hsQ15hhIRKKL+LJaqx8w4klUH4CTOqHGFlB+I0+t8mm1KAqwmRiFMbQgihWfFAyvPSu
EmPbYWsMCfjkiULN5pPYyvbHSH03QGfRNl+rs2y7UjPOjVP4H9XGZ36ojBBkT1GW6wxBchFxyCSc
S2m6k5kkEN8XnxhTjQX3wE8IITtDjZlTd5TVl7X543kf5lQO89RfZcxaoVMu1QaRDmcxxDZftj/C
nCyZ90MQbGK/u7zSooudwr7MUqZExzgGsgpiYx8fg+LWBXlaMdkSzF5qQVi3R+C1xGW3VmNLBQ9f
wrqZ+Dad6rsCukbs55I4LgpiICH3n6QbW792G4N6eCzJ4p6TepkqiTLYFgCxi6GAWzanW5NeX+rw
Js77VGW4d5hbMbdgGluXsVE+brkQHAC8unY3lY95j+VWNw5vOCZWUK7fR8KNOqJSJ/pboOjUsWdc
ZPsFYLZAr/GjCnx/kkABtRBYadGyIZA6yoEYoT5WUDG0PPSqi+BvW8F2QL2jcUcLUkPBV2rRrEzt
sIfffYaADpp4n2cVjMlbHbg6p2Sjg6aQSgEY9J35sXiMHpyhOGn/rIuoGTldlv9Ig258eNIgYIEj
jQep4MK3gnLFyVXtCgFnzMqi10z+EuxX3GQNaOT2HzHfZs0YIJTjcUlyqT0zSNcdHXkE+cm3yDoH
KGHuZbIMp8bJvaobs75RB0vycNJUc4DK3vKEGljzIDuUV64oCuOA6zrJED0zPe+/+DCJ+/VodtQj
1DElVuiyhRER/WuRQPI1nlBHVbtrRXLrHO6IMC4Gw0hGERdyC/VWmKEDGrjIUunh6eCxgMM1ixup
dp7I1fI7EsipULwgTmJpqmlkQ/sXThPHr+hFcDEXnLIBTP+jPdSScdaP13xhiy81ZnqY1PJawESn
cx6IZJbZcoI4noupae7UawDoR+pqYSaXT3R9YH4UfMjOfxHH1QshdirTG6zkKnTR+RiAyapOh0DZ
f8YP8xKzTKmzQORWHSVNW3ISH5BaWHIJ+K3ydAsgmWY0aiCooKljZbn9hCpAGEJSjVGeWJLgDtL8
CIHV5gdi1TTqZf9UW0KldUQlLm+Qzlw2hLZJvz73FQJsQOXmybsSdZWyP/8SYJqtIgRrPRKqi1oI
9S7qqXtX614Gsqzie71Ht/gaPUUDO1q9vV68KeejCuIANkFoxiYrZGBBq4r3wo8FZ8tTgsgkTKFP
5X7ibhZ7QDLkf8VJZhoiuMHKRELHgDCSxOGc9i9pvhbRhsTsbGX/q958OSJfJa0aERhGXb9glF9e
x/hMwR9gUi7RPZa5itbfALDyt3WXOIBzxpalGnC9HjVlS8qD6e05oNKEHnYAB/E8hGxfh58kS3qq
HGEWorH4Aewy7/S7yBb5gHgrpY/YCt8+oPkm4Cc6xDhthRLZbNkqJjyLlz6aCKkn/MQJyNOsRVTz
XjBQ+B/RKuGwQOjq7wzMsj+eBaoKQAE9tY5dXHHaJClwgVtDCXt/YULVDyiNCRembmEDHg4dydDc
ZSB5437cnyNajf4UpNEgnOjJUfhvZB5im99FXDZtFDx6Y2+B36w40s8EZqIqe830haHb5XGtFQrG
f7IZxj6hbkeml+pYWbjaAt5x8YxqWZhAcrdpMyCCLGrxlyvnfEqElQ53ZKU9E+/eNR35sBMOSD6R
iQ42CWYQknyfvinzCvHs5iI9vQ7/ZtFc5DJCBTHG+M4H/hdeNK8Yqg6VYrcpfbPeqEpe1L+U3iyh
wx8vJdkKIW4ouzmcvEN+j/u+YloD5Om688nf4q3MFAFSmWSXQ2h0u8wHV9xNU0ygmHOEVmDs5UL8
+ycQtTNoWiqwMwsxeDz1ywF3BpraA5Evtsz2tHpYEXHrC0Ck8Y7DUmtpsmITRhittC13OqsIl7Dv
e+phQugLIPnHDCzEE6tiq91Z+t6i2q4pfve+0JGTb1fq6e028hCNvxS9VpBBKTSIF3Oj6c3evIOa
B4KzZ04Hn5t7q12OGQ5yatUBum/b9jO8iuPRTo5zo0wpCI9okamhRL4/sU9XiWQ76rhzX34nglMt
rzfFeg8RDQMHkTq31cyiFOO9NVD935TNgN2pmIKY7TbYbjQrf7OL2w3hcQqtpvSLtLu7JvCpGkO1
ALbi9ajt9MVH/3j/LGniyvOolc5GlNt9Ufn0zhZmerMxnqGV6K3hhb6o6K0/+9M9Y7VRFAB1R129
JhaeuJPuhZbew8gmE1SoIiPRJTq4Uy7bmn5ypgyYasNB3ThPhAC+pSgEUy9mF9uXuvTz5xKwJFKT
d6o6/vRIRJu8s0bVK1g04Qpga+rPEcnwCPfjk5NrWkyeRc+7XLvpGEnqDzEmF0tFVfdUoU8D+wYS
EYfl3DoCp/g01WwuF8npGwcyk97eFDN5/Ly1HdfhK3cE2/QAW8w8FvXOlM3qvlo8myl9LvssFckz
QuPoxUUboYBmWixwjNand6Mnq3nP5/zG2gvW+rBzR6Y2RMbKnsywDMgnoek6XvcAMtgVLn58Nd19
H/kvam5rx0NwAGJRCRZmVNQRJ49Ul4Cm5dD9oMT5IzmxuvonwCwuU0QlDvpJrAZfIiEaFI1niuX8
yhCold2+Q8FtAiRoZo6LjGJA+f5T+DzOZ/BCrQ3b6vZPOLDMp5FPpbtSv1BWpCL1gjKXmVjADyVJ
XVVZ1ukDhREtkVLG1/Frq41QbIdBiTQ8+/6G69Vxiqv+fzNpRJJ72j8HH8vfFerBysamYKY74wc9
3uUI4RizQm9C7VkpDaEZDoKOKw7XdnevxrV33ucQOKUfr0i7XyKOiVgzuakPrEKLdj5fP+zPXxt/
mn3iQniscJU2Am91RRdSyUjZLFD1OQVafcQB6xq9wRd7JxYlJjXqDZSJgDY4j62hSC6qnlDmutyn
Sbr7XpGThAbucUt2XLsABdRScajg+Dc98sYdjCaIjv+9T2e76fN5CwV2FBNzHQfwGuyUp1Q4aEQu
qlqUgwdAsSEO1WrLyk62Ah6T/rArzIE6C1yOs7zLrTAd6j/YMxeljBGBEkVQVg0KhIaDN4GLjM7a
CsHebVRs/Iet8x9vtwOI+kHVqseHF8beBp6NzrLtSwiQA4p4G9dZMGBLSuoSsmU7BzQqc8Af6Poz
il5DhpSp41JEjrGVSvpuMJWZie9Ft5cqnCVJwXy4NsGaTPaOZ9sacuxlwBn4SRA8NS5XAdqJa4Wj
avQlmFN0KM5HDuZUK6U7HdnuqtrUzJXbaa/mnfihY2WLfJCohM+HEOcyS//FXh5lSuq1GfSydnYa
rrEOQ8xj0XyZwntLnSWaic7LNBz7KwFukoy2GNzMEzAtZw9aME9qrYNiFNDUX2WJdrasb1Iz5D+i
VV3EpIxt9RKX946ZmLcCw0Zm9upBNJCC5C9963HUOEDWGBaY3zxR566pbNExpLPokzQXK7PmPnJU
q+l0GNm+vQk08JpyLdHNomOKU0OPbo9OQlOSCwt2dvtpn/0rKR+vxtDBI5qNVxPbZDGqZumVWCII
rYJ+jCAyZkdlnCXSiLiNOdJ9tCe4R0NsiQHbEo6hXYTb25MHCkHGR1VvBkYnUQbPkEyKJmOsNk0Y
KnIoY9dwHal2rZuIkexQQFUZKUFBFcedo2u3uOzqWw2ebcg9IcLY1OxKZMSE1lBLnqiwWHhBQxcz
JVKzabP3Nyh4/mdYIgXMpWj4ObNpCBGfy9A7eznXRWkZ+SrJhAMZ4YgJGFqnXou1ba8chAvP01Qs
qEMVDzii9CtiVljwUJoR2W5o5JAWqnNRx1k/zNXNHkPMDT2s3mWZc/jjNJfgaf1tLvYQd307UQMr
/xgJDDq/i/vIcVB9F+ulcoCJzQAXi7Rz2taADg+qMnMcWVRgbFRzxl6kLScoCx2xBjNFMa0/Trdy
V8W6nDRJg5IFsuKnSQnJ0W9xcaqaFLOeU47o4dZk09Y8X537aJvf7ZO8NUSRBiizgbvPcqDEVVTx
Esm9N8Vgi2KqpE9jsuXPfhu3tqC5GwDqf02lr0wI7ObGdVMgC7+hgI4tvahWtX+HLKow5y+hzcbq
NczSo5ZMcoSrP3PaNYMneH2VHMlAwMIvKGGoMZef9pra4RhPpvyyMB/DMgD7pztWUvWwYL5nKhVg
a4+zEFHzfGBIj1Ib6hUmY3vOMoDIhiiFBHOrONCUveMQHHYgDJgjp/Bx4yC+ActSsMGXLICeS9no
i/KydfIbTsg8hsNXafpOfRURm2gJKJJvQjB2dOE+NGMZkXxQHxoHF+jBHDaAxDECwwin5VGb/AHl
jC1FpYk+ZJOidVPsFro6h6dNeBt8DMBveKdzSypZOP61IvdErD5YmRTNcf9IGf51PH29aPO/j1d2
TBhNStGWjChJNjiXR0YWnNOxZNzbrlHjyb2jCeX+T7Pqf4TeMJ4SlhqCZ/IcFKeGSii0kojOkY0c
VfqxhVMNR1U71soCRuDEwJ8xRbhhEaO9kpdLPFlCzUjPwJo1sA5gT6LmMCz1YFgThydECvPGDFbd
6OJvvTcOlfT4H136MFuFhYtZsTDobQ1JCgVLX4PtmbWsE+Hwk1FGV0zAFQpKQOnSLTIex/i3emtV
0NthCKkcN7Wqmro3OXd/+OIE35PFu3qmj4sSR5z47vfYBP/Ah1eTNZBbH/KOfMBGePzXLT0sF1rY
CTfSaLhWud/bY0HAdITIRWeC+uz84CUUSxM+g/pTuL/y4LZe+e7thpbJMQef79lYC8xe2dfRKKck
WDPozmK5g7CnOGhHTkWFonHIlM/TkW4pu7MGusUMfUiOmyAK2Z5EAp1UC1oHs4RAAWBKGdmQQvoU
p9wLKPHns7HLkROWyoiyQdT1IqwMYmaiQICVoeoNGj54ISl6CEwKKb9x6WBjbII02hGI0NsieZQk
vsMDvvsQEtXN5OnPBAKZ3ElIdotV2k5CWFAGXubXAap2urZL+IA6VmphcL7Ju6R9P1upUaiRsYIy
r3WCpkJUy81j9kPOZUUNiEJhlAGCwJD1jK0PwUTch2YOJOXCX9pfg9o3LL8M1hz9iSaI+IHc9rLi
eDuwHCRwU54JWTq+3yo+RHlDkFtKvdpSzoFNqe9x5PbjviRQ0V3UsDz+a9/STYq6vai/nNkM/pQU
tM+mRIyWSxzKdx74N15wTyr+gezs9rF8T15djXZ1eHYpUNbVee1F43zSedwrQSkW14IGZqV+s6Ky
ZvWn3aNpX4QkW2j5cShGynqVtYILKGwZuuKMGXqBAhGlTSedRGARA+WuoKzR4MfMTjAjqfe1hRj7
IJuWTYJqUOymuwElOi0TAYuM83fL92uxNTunvod+ITD+4UYJe18CBu4qd+RQMs7EULKvXihD7qs/
sLmR5lpUpeQHUSx/8uKyUxQsEiArjIqT5QHYBh6HYkbyNVVyAnN3I0XhRX1fz5v/iqPPAuDucMDy
wD7kDezItkaz4XNrcHbipsNgJ6YsDRalXxNJm2LxVlViS6F1eZqUqc5ggsNf2CzVBSFOlY4kP9Dg
/n3jR3xygSv2Dvf1zL9/iN5S9wq2UZzGTu9DdpY/uS4GSOT5vAMmpcj7x59CQmp0tzVKfQ1soda/
4Tmf5gtcGLRQ9rlOPz3rNuwBnrmEf14Db72e3KcA3rtMqyuwkEG+LrfvGf/cqokbdUx1ohzqHkF5
lkZ1iQrvXZlrvn6DJxjuD7PX559dAnaWD6N9245P8d85knqEpm5BCoulq1AP0CwEP4PKkW2EZ2G7
oj9djuROameVHNzZI9qt/LoDLVfBnD8C5AjNqua+JbH+3y84DY8RChGrvPNpm8ay6uwW7/e9PDN5
DjQ/Er4b4uLwW3oxI44nsr21nUG0Sa1+I7qd3MsKOF7lkaP9T93d9sfbbOJo+C7keejMw7IKIwCb
OyFY6KEnV9AB1FkRldRMEDjVzz+0v7CqC2miYmNN8o++ejuMaLo2dYTLmdq1xIUpZ18GoXSXFx3P
tZWyopvHXDt6ZBmadGvvt8LpTq8ZTbCS8wOWS00VR16FWlfsoET7dsC/376VmoLoSr4QAdflM4Dd
FNKDWMXoDCtp/6hkgbm0zxVrRH+LwTdXn8ibla1vStZ61rHzyqypKRnLHQMkkmqX8avzhceAyGyn
wqT0WJoSkDtRnROkYjQxTvQNYxMDjULTXI4uxRI3NIsAq5MZ2hKSW6RKHTHZrQsPuklodaF52E0P
RpWz3Jx4sqlmLlatbx8SkKoZJH/JQYa7t4za7JSYBG/Ec/Z9F3KH6sxVnC2pbWzdpYLK2tUYYFLS
OSgmertjZ2UJwA9s/bQPumliAK7QFSyoDwvdvgtkdtAjUzVZmu2xdVkSIAPT0EHkASCS7HuIVeRP
KuQlyFlg06sTuiuryz0GKUTElAmgA9XKI6uLdpJRvmazCZ6DskaBfROp+uC3sYJzMXLOUB1kTwBa
GOY+OZ9r3WO1IIKyI/L32AeiT6lpPJxMmBqIZ2c5s0Mh5Uw9QO0n84cPloCJL5YnSHChvSviMsmv
2JxubR0jvtu60lGlY60xy6Uj8rRqLqwRKHvDEYs5Te3CqSHIoRaRPPNmSSLvHTIHksdg3EJDKseD
x1reBRY6Ouqm4S0fiEwxx+cBJY8Rfwt+6RrZgBEamACJFiDNZ/xJTjQQ2Jnr54NKJohq/3av/U4q
frCA0dtrbiQJPZxTo06d4fOeXl43+29aK34jnlZDD44VcT9nqi4TeeYiBLGNwU0SlxV8Tm3lavoZ
nEblEKfPonyo3lYttj33nto0NKVgFSvGQMzEQBzc0i3Ku9JMYl+Jp/EKDtksxfZpL569NtEfjz6E
YlxTikZ2H6pD33SLSTkwWznJdq1ssaoyzFGxIXCDO5v3c4mjchG9f0RWTwg8TAfPgJQDD8fDyBOR
J0PuPW7IKg8SG3K5Coe4bagNZSl4nUSpp5iWks9DF4dV3XMSuhMR1iBO3iu1CV4ACn0GkQHCKkw+
CJUZA8PGXrhKJnyygAKRXTiG9RKkbqMkpgQZqdVYVgZZWbUcLbaUSoPYhzWj+5lDtnygcRD++avQ
hEN8p/ak+xitIiQIstaw8kaQBkzJ6XSPK4AxqDQXOzHe8AUwN1ccBSzjh2ErqP7+O7I4CMn2jy9i
Q+lA93A126XkMKA11YPnCGZDDMGBAwMGT9u6ezMLXmPbyk2xIZAIqvapJLaHXJ53KcVavTFmjoWm
SuAyMpWiRccIIQPBMPyplfZ68v4131zyN54CoHzyh1b+v3H0HfjMidp5kb5zO3uwstkT+v+wdKfJ
MJfeb05xB2fMsD2tk9D9FsKYzpXdLDOwpYd4Gu40f2O7Fp4BSZHzjEQkpWaloToU9fCfU+zqv8Hx
sZvEa+ED/+YUuFb79/3DPPAtB6P0Hq4IjMEuH1TOW4ImUvrgdIju4pNUpgVSQPHCo1qVzafhmJ8y
UmkbYitRblo28SNq+yWF8NI2J/DGbx82wjrmS/H4k2/OEsFSx5A/w/+5rrXp3p8g2j5cd/ox09jt
myNdAkljRkFwWIoipHJmKg4FnckMHoGjmZDoX923Ho4YLv1MxgkJr1haZLmXZup7UtKmdC2YjKz7
YTcmT7lmxjXqRd/Kvh4yErDHKBkaHidQz+LA4oHztX0hf5yUYqy5Zll8f2wq22QnWWATlXiEpKPx
fePACBsx5Cwk9RvuXvpF6kWLzPyhyQfbZGpCU33KUNyWtFh73X8NbYMkgAbr25TBkKB675TDPgGm
0u7g+mk2ErivYLZUGYxcuuQ9uIlowMEghgWa6NXlOvhF+EnJUwyoCtlLr57WgwtLZUc0PoMjeY6w
zETKXovsrA6yS5DvOybW7kjL1tDM/lqEanMFt8iKmd6H8GYuDqKrBW59KlhbZo9J+HIFlFNmk9hz
nudGTl7nw6MjEadU3vMxkb6hSFxTUCzQJeZjC8cdM9Z6imbrLl1s2Qx7ycipoR+VuDol0Xsv5Pt9
xTD7YftRDxEJsP/eAekNliN7qdxb7xFAPwcom9vHPqE5d3WOgmkHGty3WBmxbgFmj+OxBNLtuuOa
5ehmvpQDvraReAd13WXBu1igTprf7guuArZ+3nRIh+MofbZeGWacQ7/PivnMmNqu39qvDk8gWbCG
fFBJBKv3yo3UkF84QYsIFwzQ2ox7wdRoRK/0lKMDHk6EPeicbnYmsc8wSxHblqKTJaI9j5TZpjkv
DerbfnaHsLtTZtLRuktrigcY1DgvP7UTrQHjLUiLAdalPckYGLHESPSpXO8IydMGL87QkW19VK2f
HmbafWeqinjcejxYftRGXwd7eUC9IexgM3MYired0+/53wn8LUCXNZyvP4cJ+DrQi6doeLRZvEkD
nb0Xf5VJYAnH/55+7fglDJm2jkgfi5FlIy5aqfyPXjwcq51bpNDLxhG1YAylvDKd6KVfPoyFCSfP
CWQnBCDct8Q2WtO4Gho8TMMR+bZsGCrwVOtE6otC4uVOoU+JuBokx2GrDNytb9lMcQs9WP7HSNMR
wRdTRX4ZWoZXML7wHNp78ak6ob3ROpNR5a4ev4H3nmaj737wO8/DiQc0fUwbEpvjJe2l5KA7g5Mn
JQsYu3mp39ecEz0GcBfMvqo3C+eZxAKyPpJCXKYcmElqqT00LhKph6ZyZ9PSFUWBgMDqmVIxOuou
t1bhb2SWGVmjuAILuYbN36hSMSjAwcbDNV88GM3pAcOLtvSA7VUMQg1G6HJ8R4vO2c7508EP2EFp
Pb9XbakBNwSAfLHxc6lnpl+tGtlFAFsUCg770vbGHTRJlqVQwxO3ssx0DygsgqJ1s13zJ/9/lyqD
iE03YNqPmiTm282sY6lR5apreQ7FN8kdN1vi4MmrU0ktmzFyzow/ElxCVGecYQ30qGb9WkDvcKN7
6gdFs9kW1m09ioW3pxCM6X4gK/gTbZjpkz6MoR5m3e4Dwg5Ou2FOvezBdT3gz2q9ERHOw06njAjA
Xg33FjUB0WZ5S6Y7NgDLbTG/6Xk8GwURmX2Q4Li/dZVsEZKRoLFDJ3crteCcs3OVbUfoXx3i9mHi
M9Z1Z9RuQzVP5UDRziI89GsGDdlDE3XOTroehHukjop1R66H8enGCFjrrjpn109wHIoPThiiwRy0
VJMwetskD9h5CPx9iMGbZCA6tNvU7ogV7JjG7wy401qcoIeC3iiY07wq7NmaFTdmGF6jYWgq6T7O
LjQY3Q+fZS8J6uy1z+toUX1LRzfnEFjZWN0NX2VqHC1EGVVfAqaJJVJwtBB7sQbxkJxvoINaK3qt
uYXrB82X2uiWsiG84vWKuzLCfIQNcLov2trk9aItNDaFR062aDfL+6SIj5acGGPkUpgQZ9bIq9Th
u3aEXlgh1aJIN/HyLXGLIfQ6FtjCq5TfQO4k8BclW89BJ+OshZFO6P8UAohomIWnwyjyIidSK8zM
jr/BTKpJ52N7kuli+Br0yaoWx1EvKC80KXVsohh0St6p1FBGuDcoc4gTWCd7QI17YsWlTamxLLKH
5jZz5CoQMTtQ8XLx8Q7+c1Nd30PBM+4jp+TZ46nx/uC1k9B0pJxx8cDRyOEzexRgrCZCEPMWNv1W
o4PWlXfxh8BmWB8kzqWEW4e5h2y2grtRCz47CIeFONe3x/JQYmcFBsMnzUDtpbzjd8o9fqQBAJB2
1rwHPKRq/QYTUBAkm9E63BGRUaFnA6drFCxFCdXZKTtiGagwLlnLWQno2hXFs5BSdrVw61YNtEEm
9k6e+dvDlHmsW4WblTlyT504R1jJbFmUAFl2vAXHWhEZcZ5mbZkuK52bJHd0LM471aj7VNQlf8Fx
qVnDlC5q2Aj6BYGICq14N19/CpysixufxhjIBn3K1qK1ojotf2CRo40LNH4UeA4/jEB1axJjVfcn
/9hddguYuXbW5NfGg6AYwhJsveOVjexOlVCAmvPFyg+Aj9XeVHWK6ybe9FkhdI1C2A3ylnZTiTpj
MnZ3RGy2bn8NKSavGP1UstTBUUYDVl43qguF7vfeEyYifEq3gsyJVsn0DOTx+DEMqkgqQ10TbxZz
2T9ZWXlBx6Fbk7Jf1T0044NDXsbQbgjBiFwo6pX3K0Tq4SjrFPX4zEeLRGH6YTAuIzMasvRMEaq3
t016ewAr6R3TwgvGCTjjLNumSKfyorwEn/v9ngq7vHMNUXXJraT10hJTSDbxgUDS5nMn1JzBWXzP
xPFnj8es/X7N4dIohKGrg/rTwh9PdwXD00g/2763vhSL9o1rxT1OTZ4yEh+vxHuePTZsbRZmto6f
WiIyfjkFv4/bUNWubEfpP0We/inqiG8SbBy+glMVRMaYyCdySnDSXuzSAtfTI+sB70p/DBX+4Dm5
Z1zlZ9REBxDYzhTgXJXgo5QL35wwOqU2zHQd4Qd+yEqMfspe7Aofasu0WZSbLuKZdu8gh2xzzGk/
/AmOa/V27vaenzVBKmGqVcOPC/TyZTeR1++LTk3vHG/fUwhkT7hz3j4fqQPq2M4viV2xEvGwceJI
cvFaIJQJFYXD0clA9XSHSzHA6K48cEmm3W6uS77UT7d6d+2FscOB8Dob/MoecEwpmFoQlz093kaE
4aLkw4RqXZbxQjTe9TpKHliw0mXv/pom6t8bHedDmo8U+HDK8jBr4jwy0i2nIbWoV2gegIR45JZj
3e6VjFy0WW84XK4uCoLhULBZDRQDNihXf50AalG7XZ44046iKGlDfJT3v5KRvIm6phUN96oVYA3E
yCxpqA3M/A1+T23fe90RSmsaFR/28iSxb+/+7aHJ5HPY+qhuivdOLzfe0HFgkTG3Ap7z/uUwja12
vzdLjFeGEOVnt9DJHPS2U11LCyM0vkuySZxBb8kK98QMHOTf59DEJD+k/5aZ+z6cQ4VmueIGj3O1
MXGlAGC//HORwnXUWWi4bvH++3Grav8KDKzCwweNsRSFd3xihOio/IiyhFqv2QEyStoEt5NX+Qxy
S+8KjtAj8K6VaGCsmIpJL2t+3F3v/f3RxHFJRPQ7Gh42Mjakzj8U8LmeA7B7QCJGEImlphk7F9RJ
bpEABYxzvXFsOpYTDXIle3EM7683/w4Iy666JNrVpqgywilcmsOQD43fQPXGtUkofFjDF4LnrY2l
rVVhM7G7MrCTKNdH9QY9/BNtWTfn/1Rz+I26l05tFzoGPGGMFOu9q5YIT4GROTnQYevvXj0KXUk1
pEOmQDTPF3COf/GwxlS4R12JQdMHEmGeF6YMSMGHPGPElmCdhWupNG4eHmXxnG+D6bIdkdzL3rfc
gz6VEBQkAlDlYRw35KRrKSjKhdOSQaHGvraER5BuYCpzAM/nH/3hy5zuwI2Ij4uDHZX00yuEdjc/
UfX2WvBmIzmdHawuAv4d4/Vl9kyLDx8aTbmfch0iEtAMsn3Yg145yBE7/gb2HRDvb//lEW+vK+Gk
eO8KrSgs/pUzJdHWtfsbcloRjt+dcZd7TKGH6jnprXtdq0xP6u7SZfym0ROsLxaVP77c0wfQbEbc
YslX4DWIttUTPMWe97S/qdJj4P2/EODSisUsZXrd9N6Jg5/NvZS3DyKmsG+Y+zuFiIrmc2gsjYQs
2HhuBkiFEpOEvjZtiROW6i3a/S0jjiEDPB4Krd0N4jfl+m2sgYuty9+Gha8w+LEkBAD1CwHSqIOX
9acaIUqgsQJ+3uHktNsRBnjeU/8K9CcOOBbU0fBe/rLjcDjLUF4tCexxpXty9v2dPc4KwdyQAGrN
Gyq9NHH95Q5tYYgjkWhtUrHQ8ANW58amWHUH2EOT8bksMPoN6aDkzDM5D95xgMBdrO48AiqBdgiH
e1e659j2HJv6r7y4YQ2j1Uhu0mBuzA9Sfs/ReRx2zpXmC5EoszkszRncOT+aK3sChrEB7ay3tBdn
R+riFKBIs8P/SdrUg73hHN+Ok7EwiCmTUbREc7JbZpuKfD2X+qSIYAnxGI6nGA7xgsNv2KMu1xTD
BLSubJC0GYmc+XPIj+4sdEetE3ZpeHk/lFLIzkHtVo1DaAjugClkPqcHoIhS27Zw8OuZCI4wQ0KM
8PhW0g0S2ooKbqbgAwMe39dKTVpxhJ9Q0T46DB+Lamwb4VbWh0L+SQCb1fF6HTXuy3501XToe1yq
OtvMxp273MVuW4kKqcqR//VfFbYdqDoXei7kZjeVFBQI1rPxmDr0Dgy+8QeJUXiEtfEqpPsoYiZX
thG4fg0Or4HLbOhwj631LNhRBPZUVMvhWqrNFO3Qzi2mPMoFdOok2Vd60TLhI8balqVYNPhHIDJr
hQNwgshBmulldkdsj2hDSxs3g6eBoA8D4vNmghDGOVjeIfqSF6YKq9rKplodC6Gfzlg2cROSaRkE
XOELOhITmodLPClmUUPF6A5kYD0u2XbngK0OdDfY1CVfwC8Fw8RP/J7AhozBcSpeQA+hPG9UL4sR
4i5vIaNm7kbD2yH586jvvPGe+Gwc0LerW6HQRvfTTsds+UlmGR3RDfr1pBd3avJwqP8Ue57rFK+9
IaNqbHivsDdoVab8f3D0EVDNwBgr8vd3XUsAp9XStfdBedErTSawEXMQCXYSN11HpOSkbmX6Iqfm
T8T4fHGFA3FpHUExuAhV2GhZmCegwxe0rDU9fozLZkpj6xPJCvajs5p1jvuyrXs+Tri+Kf7dnInF
62ABjsZuo0IQFG6JQ8CGh/S7ltMx+ciPeOz5/5hSHCa4U343t1rBFQUd6x8pl5227X/Nkwp3Lwxh
xyWtUJYbOOYRuN1ESIamT+4GoOmKY9+3R147PJfJ2Qwtmg2Y542HKi+ySTZBTaytR21GbR9EAmZu
ugmZWRShz2b4SyWOfLiH4rhBwOOs9xT9pOyPLoNdotUuJtP9Nlf5M0MAM0PtqsUD/oxaOj4KcDrl
eCjuVbO4g8HUT+ReP/cGWoWxP9gpOJG80prFoF7GrzPPhL1SMHxEOsNRkc3ZMyAruKr0nxeFBCMN
xFXj//nb8Y1Bb34a7pelDXYR6uH1kB1FhyJqwcpzQ+UBpVHOnpaKBM1axVAyxWLLlE4tRHy68/ut
aaJzOJhmdB4GyWHNd0GY6LsdRd7FNSJAaVb4QonzeA1a6ZtjUUpojb4s+NOaIvRBQDfvmreEgKKY
9lG0A5W0/KCNwroXSd84nuUajb4Rxk+LnxJSDneKyAaWeIDLWH4CICPUhMAVD0GsB70y9EpQFzSv
FuKVIMrVJVjItjCzY7XmqMwoAFQGUlQ5qPfJ4AzjHufXKICCw/lPQXBIKsXhFAJLATxNy+/iwdVH
UpyoYKrmvMdAGOS3WbtmbKVEXYWeaU8+mXZRTeAu891p+Ar1lpf56bXMdVBznqt2BBecAVMHXugG
mtj+wnr+lsmihB7TDcjYGxZWF5T+dyAG9XXpS1uxslU9l1i7OzcXGmjGwpDv4fI4pKJyBgrwczBZ
Bhzu2+DYhluZj/xB/Xjwvb/JLe4ZeM+h8is10at/A/RUWJdZRq5N5lbrOlC4/Iac1nL+NYaizrZS
P5w7Cfz7bpTg8Ghrov6yITrTy0CSvUTf1u/B2CLWb56nbHgj4Pzb4G3gu9RDHIh2R+hz/6XJV637
D0MIrRWniMqLB07uoxQLrA4dsQYF866LJV2gud8BoqyQqqY2p67bpfJ8g6EXCP6Qr928XroQSINT
p6RBcsHP3DzSIkvGAaewfuRHMHvb355T6WESdJaJNsGdXYAgnl0/ZCRCQIzYoynzwczZFiLru5n0
xBl89uyCfKcPtGUEE7f4s22dafwJw3L83aTJCKBQoclVpJqXsTpBQMW0IkgGxJ56VSpnD93ni/Q8
Lyyreej9rT3R8Vo5JbhwvFcPMxV6Cl3dm+Q4UhTEJNLXrawmAT6SuDXXf+4QhfWuRz543Vs80Y4/
cMh92aqV85BbxwiE2/oCGukvfLa/BgQIjbpFwLH2LyORbuUOkY/LJBEvpANTYCU7ElJTJaFxNcQp
P5Xxc/FHu0C0CPKBmttFUM8EVCKPX1FsH6Ahvz6OpGTr6T2UhWD4UG++rr36YoPFt4ELpHffe0qG
qP2sR3VEXJ1zIgQKmIiMxNM+uOaaVhNS8N/TDEJQe5jJTuIBGEDLxxX9YRbWqjEced6Wmj1v0B4O
Gh/2dXpJ5aKTgkv3Na1b4e+FhzKdM/oIj8B/8K+/AVuFqWYqA+SrYn4i3bVXc+GynSp+b4kYjMiD
DNPWjam/aePTnyGNNY2eVDJxjVLUdbSFYFiAMIQQ5b3Um2kxljLHoSkezMHU/jWx0Udzdc0lWr0Z
eA8xxuh+w8GmFF3XulQqC/9tioM51UY1Fl5CRju/8GmZSt3gZgBj9JqT3ugFwn3BhmDXov2433lh
b2jY5XkwaGGN4uxsMn9hcpXru7c3nmvbAPI7I0ccNYEdb2FejNq48EvJ8Ftdq5jpt4W/sN0JeTox
26HrU7XWpHvosESk2ETuWMndwKASeQ1/LMfoe9ZC84B8PDerIvVUB5ljMQk60txv2XV22P6BK3kg
1FjIfxqWi9YTB1UYLGNSWMKfovq9QkxJPiC+Uasukv5/xhmMIh9kzswxxsWdqUo/ZW9ismNZuKLy
irKlmb/e9zlliHAYZGHDUAjOPnUIHWEfF84dt1debBSqH4pU29zjPZiXzD/tRkAaLoTgt0zVSbhd
eFYwHUvyqHQTWmBQeCiEKgsvlAny+iaYklJGez6YN3/9M60FUMOGzp+teePeZymrh90j9Z153Yt7
4Juvp2KhaVdwhP3kuAT8octJoKCFiVtGAlYwmVhZm0QDL82toJgMaT7WsedhfEEaqAXLHyLog8h2
/yK0Jk6MuGw6UMlLxxqoJy2GP7cJUwgaH0Nvgqfp2wadkuQEY0j3Dlik4+B1rjz/n0VH9FXQrQ1L
ScLUTuPWsgTGM3FiMdNs8ebh1ZzYKUdOh+MRmVM/i2c/r5fV+Q7e0SP8MlE6LHvLw3i+oKagyrAu
lrWRx7IHAOc05YmGAOCXp2p8YLXR6IqbtU110pWR5m7QQYSvH4oj6E/d5fcOVWEn5BzslJngdQpf
kDZGXrqI8y5+7atEiKqLpOlBfI4CbNpDikcQeEHqz6XAfizUvCbAo+HDPWnTbGceqjBVbbTWnVY5
9QbXx9zhe85UBjAA3Uub2eVHB6KvdmhCH6otRnVNA6GoaGBBoTRN9ZqXNJi+i+Xui3PVzdzyEdCg
z62kE7xidA2DiA6qgQwzPymhQG+Idtma806J/8rK0QgCGBu6l0hPvfLztebg3GzlrhSjO9Xu+X2h
KgHY26f4lzrMIMx8HJm2NvVWneliSS6uMZO+ROdD9GzjNOabhbPb7m/bcbqcqKViby+wnn3uXv1S
ZPibJlszCTIcqCv3yWeh19lhfkFENCoMpvADNaDdXU36K7xjpb+d3PV8Gi845ali34MubTeNMupR
8kLWL65zdenEPxl550RY9jeCXpewnZ82doyjT9kFj5/aJJ6SWfGURHIIUeUJHanm3me9sQG4GyFt
Tvlip2wkarl1a6NuOoYVk8JjMmg4AJ41sfU7jqkholM0LfV7bPV1Gp7VpEWgrlFQmYxGCaA6kK2+
tIdmKYn74YWE4zZOomLeEjjsS5Gek3vg5oEWPjWkUmoc0+ocoAhx6h1jSI/gVrOLq/OKgmnyHroq
rMwEKnMlrVICBi+v/T+5RU1ZYN6unKJJjfHuYvutvaCWSZ9XeukXQGEXLGSqrtLE0oKp6PxVt56b
Rh0dyl5cdBeEyAPOdZv/lpaS8NkiS0GjIPfmlaUUcuXw3JAzDkZZ9lUra2kikpPjoQ4Sz6L0OJ1N
Vp1F/aBZ5UVZpSCwQI8X/3wQOOv2lbMNHt2obclJ6Dya9pZCTrtw7SuKkfmS4Ntftb4CxEPUiNWh
LNYSun0q+PmNh/blv3OdsIxErmF5+uNmPvuTHljDmilgVC42yLo0OZqvuJyihri9sWAGcdDc5Jcf
zRotfWOl42Hs3Kv5E1c0vV2RuXZsbogDqZF3nPxQFeTLIbtkvlzk6rVVwGRdqKhezBpyRo/JPqwg
EymuMXYxeHHBEVvN+rWpnVoMvft1yENhj/AVL94fUHiDxT9GvxDEAZkAAOVe4JHDv4tcxDIFBUZD
I39pzOoUzYhit0YzvGYOu+mz7P6fKk623Z7L+PyVFpmHenyVRWJX5GHhSc6YgYMiOCGLP2xzlwYV
k+suxFAbZ1Pzb4Bk3ojr9ka51o5Lia8x1dEwAsxd8ZFlqRBtPhzlWcWbSfiABsDtB8ZW0Vm6LGIy
8iQtX6XplZxeZ5SJevlCAl6s8X+GzmZsAXIRhHTpvgfX0U6j7SitUFrAMuvd574wE5YaMBaAt0Ad
Z9wfLG2l+3T+dQAXj2d+NlLAXPGmyHd61sibenT4pu0bEYn0OXLg8Uoli7fLdAf5DljKpQzrgmjP
XKIPQ3hDgtqRdXcR7N6kaLgbFMETymoinAx1AssIA7zjjHlIo/fFge5g97KO04wPnuHuRX74+Ol0
vAMDaQv1bHJzjOMzcsrV/F+QY5leShrZfSmicWN3rFQ3Ct3OaXuh6kJxc9d/zThskA7+gMQoQ7J6
XaBjKUa5TdZrxtN/J21FKTPqxUcun6p3TiRobVvoG2BgNfwutKDNyPGNpkD5X0S1PYqyGc58+0+2
MGwk//bLABv8ET0P85lJr+KFhMql3zvXveO/OXgQDd58ypOcwu9JCcK/aCJRGSlxW1s/x49OHaS+
NHfAtcd0xKxwEJSK/A1DeQV1yBQz0YgQ4dG36wDSVMbrqtoYhBd4cA/hQ7P8/+7RimkBNDnLL00y
3U/WsSka7m1Q/3D460sr874AjWIsfYl2B5PUBtSPvADr5gOhYpb03XTXsSa4BK1PpZk6v+ozEKc/
gdBI9Or39KbI6FWK2w/Noh1LtAA2P9Fr4MVR/2dalCCCkYdvPiuU5PI/Pipq+uWZj8L+tOsPHihN
4neEhUV+J4/mm8efrw3sx60jHFdHcHAC6FTrWQ0N6XoZOgi9xfi9Z2MpC5YsZVZXVKttGQDZHxIk
lDOXY92p+0akAlMcATGmlqiPke75NWROgvGXO7tVfTKm47bmcSg8/Zp4jzX7OcgOm0CxZay1pTuM
odPmGX6rOrZWxAQRjr/RmFh4eiq6Mi9uEO/E8Ywn3xAODy6QEy9efX9EdmTkRNr5nCMz/HQAF8RR
4fq1eM4xYKS9NyOEbH4+ta5SFl3Y8lUXaZKqob2aH1txc+VqLuumpC6R2u5jmpojx3obRWhlO9U5
Fj6OMrxhi2Hn31kfJPPHR2BPofQi5faxXRVENMGq3Fng/WsqJvJ2pwxGRCJKYLmKGZQQUXGe6ses
7/Kd6/AkunqDcW/TPDJGrj3HZY6SLeDVsndN61cScCkcNoxGiQNx9DjkswZcbKEul3z/Iz5W2p0b
Rorqz3mYc/tFm4/k6x13ZYfDGYW6iyfSl2INNGiD+HS/SnFW2A9bbte5AMk0bQ+BoHYBSynN+tlB
bN1yNTKfVwfLd8WzTaWBZ7WAA64H6Na2tiOlX1pjT7azmvb0CsXUP1SUU6q9lhchn+uTrrfCn8mG
c31OsaRgmxs4/pGguA6KLqc6lFO3ClgLQHhqv33KM5mWZjqwQyGoxDH2xLsqcvr4zg2Kj96VooRi
qYBOsHJcN1XF4tW8X/lidlSOMibZfC6ZHluttzg7/yj4tJWCPq69pvMw0fNiqjlOjrA31eM4wXa+
ZSTvbQ1H8B4Xq57/9RqYuWQGfMEiST8Tgj0IMd7HKKJKRzrLuisggIdDPG91uR9WomyNYq3djdHT
3lrkzE3FBYaoDFTkh/v3MsOR0sPPMydZks9MYpZcBsutbuM525wmt3r/febeW1GI6qpx4Z7rUyYR
6ZpGfkgZJBBsWzD0MX4fkMt6nMG6JNp+rXSchwdBTM02gKp3svHn7wvf8twll5LqECFCOnP+tmq0
ArX1UfoZMI+fFJDJM8jMndQWezfYo+aZJGkNNGkzKFS8H0jpArsZxx8gmkTW6jScNej4/ONhnbca
oDn5Xbe/lB/65LASuxDSdF4hVzQiZn+SdvgT7O4IAOtkC/yJ9VfEwk+J7cTiZDyKTcv/ds7SFyJB
DU3Sy58Zj3bwjpCtqVRtdNAaLHT8h+//hY59BYNIkFNDiASLWRX8sG/GnY+5gXMtcDyNPBZ4ek+Y
bErA32zATaU2ZKk3UvNWs0EKdbNaJ5iSE0RpcaxCgJ0dt3glMaL4HTpYJqbK7CCn73GFwl/v/iY6
9VLQIvCczgzYBxJjk4zx4xHf1nN7fNJT0vy/t0vVToWVYVeLGPsj0K+huZGPT5keY7dRkigJpDyj
g4CnFr2JFVR6V2i0N9LgzlPa1m8IrY+Sd8W2P7OFxp36CGIFG/xlV9oOFDYXoh5ctlsQ4UbnsjAx
l1q6clW6prkv2C5LO0ISpvJHeOMLlQ0Lxk68YTOFtPlqe+IPsjlLEKy8ISy0rNGngnTfEdegQMvL
nV9zpdhMD6DcKoMX75GC7JwoQBLH++4Zs6ZnPZmd9Fvi5JdHIu0XoJEnl4/Cr2LeZcGJ9puXkCjF
YKgN855E9/CSukqhslx+6K6yUFY/0519QbSzmC4OrS8x5yEwsh0JzXsxIdGxH577j2ojzCnYD7YK
2rGvXSapHbiv3tqjLTjgfV4H7zI+pWZIG/L59BD615jqrruxnCrKOLHxpZ1DUJ7hzNRD+DQHaBIe
HcyQ2iTUliGe/H8MypGV5LjOJXrSyZJeUPBDiaXoVWbxfc3XolXMEewuMwQpJ/iHkpkoPkExLxOk
tTJvZXK0o05EKtEoL4BOSPwOvgzGPmSBtEcnQhf1pwCgGnCrBcoRefKEvXoliDryoZnpMQlpzpkW
rdAdkW6p4nv+thQ9TIApz/spBZjQMTiXuo5GwnVVGUs+dDdC6/JRQW0WeohT6nm1Y2WY6EaFelRn
ohCHivZQOf2mB9x8sQuDlhuPN8mtA+XLIQvxqtGIamPK6Lr5UWirwFbur5U3CseX9Ef3x2HI/eht
sghqqMAJtUSA2/Y0l/XHyKHPYOdi3OZy1QjnHuLmnbU1b8I4Ty+sckL/ujXbDK92rBnuNNQ8vOdk
kxTsAUxKIBOydTZPsLONadexT0zKnV2738hGK5gKYlRJyZj6MoFh7MvmQ9gFO1paehi0Csl2wfrI
4tBKsw7DahPzD1hQpDQkJaKGmj4dtifSa21DspJOeg3JdKSRoUrfHqBwXcsAnmoFnWG3dRvyBnYY
vCmx6gzH3zjiCVgAylqyG9NOlI3aiXR2l9S6+6pg0j6DaBwoGJhgHyA8LDI2ImO1wnwPLY3lF9m6
xuuTer0E41m9GhSEfQjT9+X1EeRknrgIET+kFaND+uEWUeIYXsOtnBo/RulhIgt1N8DxLU9Pebq2
K2QWPb73ezsgpz2gINmKaubcQk3x72/KNeWiwSvfqFj+6HLer0mGYPlnVIrsWnlRQgVtJgaoeWY9
VJ4zCyEqHJ4iSmcpGiy3eNhGByVvD2PlcnD0eDK7Brp2GZOgcgKnRiU7ycXnQp29P7iGIueUf40c
lM9+yWvPvg1TzNaR7jHcmTL7xxuGgjc9tAn0qWjD0TTXtupW1ihX0mxoj39xiu8hgyFl740f0hMO
BmPWHpF0o1O0HGTwbKMWcIt++RP2yPqM2WZe2DwYQA4hKuAy0deltXjKgrsPfiOlkTCbS5VUpKuJ
SS71aI8wnokmvvWvlEilWAGDYdwOiBncEoxrh0BveflYuWi7fW79I3hEcTkNvEYJc5DNUCgK/Pee
W2/KhpY0dpK2iTTXtO9r5UBVI1pRtGWBufCrOI3jFXoQCr5GdCaAbyu3A1/BYNOyyRafjIGxIGVw
SfEFA288TzVWb6+cutp69StWA2ZzsGt9dXGkkYZVKsXOmVkmQfXxnNGXxjKfsfMySH532G18VUz4
uXlrm1WXIWFTrvAmMOgfsakVWaDzn5bW5kHd6qu25A6SCimo4P5d3RN3oI5FCQaaDVzL/Rm5ZtHs
z1M55hNjv5bnfxorR1VxreOtvzLOSwKU30LkMa67rkTu2nAtEb57jC1gu43+gP1h9cytyzlj54YG
Ta9NNZR3mqhI6qQMd78GZlSmslDvpOnn38RCwxKIFqzbEZKEh6zV1sH1/nhhVteCZsa+LarG7V0r
vLGppc9Q6hxA5GyoGM1nJw04DavXHUpoI5T80z4P9PQ9fr7MxTbVylstlQeD66wRHNc7VzA8/6VI
qjnCShjHtVKxnZ76i5egmicgdDHTznGkjYMNrI3lbrqLl8as2Vz3dpWNjwcnUceiEgWDX2dHNbHH
VxLl7gff9kQyE42CApar2L2mRjhHrMiyw6kQzQCoZOdE7Mi6/WRkqwWMyDdRdCkzjvOK6j9V53C1
VU4XFSe7I5MA+Xva2zGxLNL6KnemmUFKY+py+nD0jv3IkdFx9MO3Hkhnl1D3T0ls7HroLhG4kutr
kB79GrE59UZceotW0hnAhKeBZ/cK+Xpfy4ATzNQfHs37x0gnqlK2+ovFuaOu1cQKHV7Xl3n9vn3N
ruAYQzInk/ukq+/OEVloIw6ID1OtZckhgRrO1p3SDsxR6OhT/lqSFldlSARTj3/WBfMZoeWgZ66n
1d6/5qK/3ESI6Qelg0iXT4tH3VSNvelxj+ZzqA37JnCY2B1VhXvKgutO1SEKeQEM0KSPf0vpM5gp
U6piDKABgM8XDHJVkRNlwMB7Cdr+fCc+cazSJ4tkDxFy6826v3oBkAApSXtiZWc5/j7w6ObVzV2f
Jgw8Ljmq3HRinDPCChQ8VW5BydYjVyPYu7GuyRYQcK1wB066oYPC1ZTw5z3SFvf7iCxoKrOHCphG
SAJlP4OwTMPQdS6Ugv0XMN/Vs7Y1/10sxJHh8B48iwty3yd9jY8jCsSA8TUmz5eFnu5SZ9aKsOaz
xkThd0xgWhoULEYotrkJ8GjdP7B3wgs8Hk0lcX1SM9dA7k1qUlmu2rh9INVv2pAY91SmTtyiXlXR
dkfY3ZK+69x0k5cF1jMmH5FhlWvjVp+f58DnBlewEwyX/PBMSdz1rWnnfXT3Hwy0+Sa1YH7kOSL+
yM1SQ1qMFUkMqaMFwFFm4M+wAnCwUTYRUgSItWLQuNk1N0eopKKkpVTaaWxs4tiX08bM1ttUbM6D
9WTGIoCALjIPU/umlDWbW/dajLKR4dDcvbvwANFonDvsR+lxqFvSMhxrwB3X/lYuKKq+ySbN8R1p
eBSEFZJKnVx3OUbLqUy9STvrXNVfeT7PyuwDc6iJqqNGjagy/q5cNDg4N5TDJjr80lD5wp8iPWgm
+NJ0q0Dc74QEwYCA+VSAjB46Vkzn8Kdbr/2tlXU6X1NGexeAGEu8SIxfb8Ud8R6TsYT5vgp8TRoQ
JYITSDrXiy9ngBUgZJP6R+yFNNP5AtWPv0QG5zbl4GS0Xc/FI5htbrI/9fj0U3uWZWmSWE2uCWW1
Dn1agOleQcAjRihLJKMifnP6lCTBSQwqDKYOoZXuL6GczwNtlQlHpqv8PtFrETXGenypKXHsom9j
4N17Js3Jo7rt516K2YETjsVR93zjUbKOZlgx3n6Sr39UD+WxHelB0Iu7wJWuu4s6PbJSZgzqK5I0
pHuiIhHP5vxyxSPotaijs9BEljvUJtjKg/T97wZ1IJKoHCnVkJp81lnH9srPfEM0dmaIQZ+r55yb
wVtnD30++dknksY26j4m+jJ9TYConYROPKAtx2WdZq7uye0cPO0Axs53Yea+TeCP22P0SH5kO9n8
j2z6NPVyZcPmaQ20Kmmb8rNn51QgTV44easH+xrDZStfBsn243xTqTgax3jquFIqUXp0HlgaWx97
t76CNXg0AR336ihx07PZjxwc2mnrwD/hSY9nnaErBRoHBacooOLDBqjlKPuQgv0520KqrWSzZEhQ
fUEcWdkKs/JI6hJUJkFPqtf74EL0u2I+AEPb4CxfdPVTO2B5ByfWS1JuPL7UOEjRfSS97nxkKDV7
o8/TPENIzTxDie8Q1DKpVRbuTLJJnig7BAYjsl1WVXEHd2GiF+d4C/cxl/PIA9idQgAtbfOrvHIe
mpHgIj6x9Emcs8sAB6r+MQ5O2u6p/vZLDx+eeEg7sKpA82KEfvWbpfJ0eo/NABKQxoAz2ffG9/hF
GLBdBvfz6K6wtdjR9iu/6i31SBDlmUfC0xgKarYwcJmkx4xBm7fCztqzAx5c1kYsyJ2oQtCGRIQG
vzelGo72X31tiI4QiusjoLnWaAYSZVRGY3kOdVnwuNKyUa3E7OeSxEkAqTmdBO5tDEnGUmZSXo+c
OHcY6fQOhWBitOlS3T4KBYfy9e4QC/y626i+YcmbH790kjPgeZExdfhZkcdL5J6xduBH3TBdjDCG
+vThGXaK4vLBLAJfAx8gZLOkCFT/oui/OwFoq6AaKrRwMUgHa2HcmI4R4R1dZQ2EHHMc/sAEyonQ
vl747aU5XapCKI+qHRyGwIuE562f82MP0FQSbyo8Gr6yji/WRiLtJdPusR7hI2V2e6SBog2Bs944
2N63fQKuOntGoznYmxUdvLasgmaztGqmjg3lreBtjQEgca7UxyNCXV881kxizQc37IsEz7LRWXv7
EZd09NDAIbqgGX+Wnd5Hpm7cBk2AMnUMeRf8LMrZb9/T8fc/djPP5qEkapywh6IJxoBFw2meg98d
ULa1bzsPPijm+D6X1sVgIn2MC+vq2ZzlJwpnQAcfZo+L7EG3NdymB9A/I2JEtVexGqUb8bVi0aa8
3LFMuKr04OdL8Ereyk9Gs10HC1SAct5DL7NUZQE8PUTFIWxXwcA/8mNeQXkK0yDzeTYQ0eu4xEqJ
BCNkkOeUoxT6a04UB4ZCajYg7mz6U7xJchUseSZBHeBPlU9YymN0jD4GB23IHBL7/KQS/5D17A/l
Ij1vscgLScm5HLvXy6Z6VOHUYzxR4kWAqGRH3ubpVD2ySHF1QvfutgtDfvLIj4EfSkJLcJsNufdn
eJmL7qGnMyZgsFb2UrdPp62BpF8t+rQPizF/zwVuZOk9x/GhFxHsv6zCM0OYr5aOqbzFtxlAAk6S
FltV6pVP1LavlL3a4bdTf48ulpvbEqtnHxBg1CsJMo2bt3pyPJcYTlhuxRsW6ECiSonY2XnWqN4f
M17bhrO4suomF+58mNoVRgQ7ASpEdv4iJQS13JmQeMVQt5pWHQtg5IOYkwCqzr+JXYRnykhz9ftA
VMuZLIDPNg+PS9IhtMsVxTKmh9i8/dFMcq+wim2xe0snt6ZXyK1yLssRQjIX8t1ONG2yFhju0ghu
OSALOiIY6Fgm5gcpXCgJbkj99kifdvnyvoDgw7SSfaU8VAfFdCOv389whu8ehYX/6/Jq35VFQtY+
ScFGb/DkD0mvpAd6ehXuj/60KnBo1aj6WvQYs2ssNC3o9JurUHFbaOurk07NXaIvSpHFnM+wuWfM
rUZdaLLjG0gxYSLqMhcR+mfgfJa7GmF9+dyolgpGHtbvnzC0OZT9B5bJlvJNtd8CtdQuXm7dXRwu
QS31Ac4JOVCjzHNi0lo+F+bbFGlhmWjQApkfJib1OEq4dtukKH8jRYGT+8yj8fh1zdxQLGN4uvGU
iyImRymZQInG7MxhX8IA54YzbUa4xV/Rlz6si7HxF+7iHmPxailFXI78Mzrc99JQHrWKp/Gn8v1x
jytgFpVa3cKonieoRs6MbbDP7Po5H5tZ5Ofif3FHWE/DtRjxnESJeCVEHvfbOLRhdDsGRzau5wAZ
hgrdosnzCq9Qz0H5GEjIdoHOqD7KQ/jsVLJQdojzu/pv96FBWqPzWY7oH6NuvYUIbsifZJIJEGd4
3dfMsoHD0BQKAMHhTs5WY5+KeObRIYZRtDqCWqVb+OHwf3uKV5iqJIm1P9nDF2+frctwjpCUSTfD
ooQ7kUo+4CjnxvUdlBqsIBEaBBxmShb3orBhuuN/5axj7vlOfmNcAFt8BhhJzDRervQOTD2WZR2H
ym8HmBIXKCeDcb/zE8CH0V98q2+Z5Ny6P7OgZTVfgC/DW15yhgEbPbg5fJVEFXgU2ahq3PzVM8nm
bq28n46EJNFAyp6lVUk4b3S7VfFbDSgp00w+XNo9XCm1Zao0dBlI14eRXtlVH5fpIr6UnAXudZYA
nvc26YOgTYBcxumTAQ12DhxQPl0cAq2byxtg5MR3/RAbzREqwDBA/OpV1/iM+EG77ZiBC8h+M3Dc
lBuwA6sfoa2kNdpqARpT2dg5BDAc4txb3F9icyByPo+gFgTFtXNTnM0IBylmVL/+nyT0s/PiiHHM
g0kOzuWE/5CeuVqTpDkJvbNIZxUfnjLzHwTyV6++GDIUCfuNtUcnbaH3FSIGZHJsOtg+vGHrpN3d
+CRxZGSfdPPvtbRDnQNq0sawNk/ReW+F3tRS5ZAkR8qxYDEXiZPOZgaZGpNmQ4pKUN66qeqx1UVT
a590B+qGFpefRbsfTnmCgoNKAiEKqz1wS4QJnFQkCDaCv1FG9VvizCDjfGNDxj4kw2AwiTgk+61A
yByIPE/oUwUOSu44nLub03bhg4cF3uPllKod+Ie/w6E988Nf31ZrUezdmdW6mdowFyUp7wCYMY77
p852F/TefRnUXcC0sSEcbIaQdGjepHJCwJ31ZzJ4PlH8i9CrCgikygdwp7Y8ZOGHPbS9odQTzzBQ
vMAr9CHrG3/oSuO9qYGguAZU7ImLldlzPPQxHtiCvC6ZwMuVEvLP6HLIr1yribLYMsw8IxwdjF4B
qXqpO6ZOJOrD/i/u8pmamh6NdRPdTf20t8+0cnSeq0vaQlGwhxLx7E/Arw8yvFUNhromYXuEIbHu
r/Rd5F51U/ZJGRzCrqFoOZ3sdjhmd7XNceJ6D6+e2DSil6Ozri9CVQB7T8tw5fb/4tdINTcIpp+p
lVJZKsqGytQLxvQcYv3m55hLypvq0aiEUmsQUNt6VrM37+zOp8Bt1ciA0xSONig8pTg3wceRdwyP
LyjfWtKKm02thdVGS891EZGWtOoTvPy6Cgb4ofEKQ67nH+JK9Ll+WhwIj9siOCWXF9frGl1hUrw5
jLzKdUJ7r9OC/CuzF97V/y+SSKXQYq6h/64ZrAfEWl/iPf3J+/gsgf63Sc+b2nYRoDZ6tz/bbOvn
CpDJocomzo5xYIkd+DPHPsj8SnK2ip+5W2RbBbsjuno7xbHkCAXkJWuTtaCcI0/fngmNpXRcIuBg
3t6LbmW2kjBJ+ykGcd4apHukdDWmbCuEYw+h6uLR8Ag4+K6030cQBjgN+0+zVMrDNXrWWg81aKZK
bSa6hMY3IwdtXejMtxcVYTvzHROAZ2Kjm3IaYnrECc54l7iWn63AYKUqNn4uD/PMRlPNBraHXP1B
vZ0/gq1R6omEiMStIdi3nu+D/mEmWHWSnWzEr0j5gp7MfIxU9MgIWB9gCMQuEY684Gajr3Mqa169
nl7tO31BWrgzxwu0iiw9YisgtiB9kALESdLXzcLu37c6ntk/ThZRFF08dkvZvPY+Dhmp46zAdytL
52ugIYS7AURLS+r+elJVW7LI2slsMoQroBV8akczIIs7oduad6u9VXYaaA8oKNGjaVC9uOSvRWap
ZwBFgITcF8Nqv+/Mm9lc1F9KCQ9v3sSJgCDrj56ibcDvUi7qgnsGfWZcmqDXYLbiaxVdx7uQuE/A
HelTYb0hUDosGKT/XjtuIGfejQ0oavlepXKz1WnRNt4JeBHnlT9lzGeofPBrAR5qFNzka0fm6f5O
Gr/1V+IHoMrwWqAQiyy4kXhA3FLJLABDpKoYGK1wqiMi+B374ReXAYG/1E3KiXwplmsjNAXPxUwu
Uh64UquwucUzpxDOtfWQgpap+m1wtpEpLTWDoO5DCsPUWFrZrmD+R4RXbTMphFpJs28YfI25hj/h
8rQXBqwmvNz7sm9JLd9+nNaP9nBULzUUBu3dGfVhr4EuGV5nmHgAq1iFHKwFAdraJJCP0n6JfGp8
yw+9nZW8nkP65xe1wyZaCevmf0LKDk3/ymgpCtwtKnzpNhTvfoKqp3gRKASHSRAWJxTVjzAuvBqo
8V9yflDBqxpEZlPasKNKCVjh/2uEY6O2JF2wvYoLWaJ13Iec9q9EkQPJYr3Aox/UUBe90EOL60up
aKLjy1gI73P8g1hh1up7f23UTVR7mHpFurh7QAPc8gVsfNXiVBs3LWyrRt0EEr4c5VCQXScZiRyr
22yy+HnW4n1dbzr5II9Fzm38oE1zrBi5Ithq1lUIIcqsCoUTR98jKqGA4OpCwwLye9GmKn2KGfo6
i4fOeoVum4B5H6sWs8lu1b3TS0FfPVy1Q1XklggQgl4YPr+uv5ggEGveU1GHcVX7DT4URGKJsC2O
gbNzSoheleugTFccOrjBvkwJ4uaoNl0LKBPena25ZvmjtxhrKnrfQy4OyWhW6fkzixT+Cwdpyv7d
8lZZXXbElaG57q6ygwH54TmXEsm9tk6F3uOiCFPMO5iYWraztmTd/eRzNaOF/scAHVvRzU76iELg
h2ycPoYuoc1jCoe+KQFQTG+CHuGOS1WeEmn/IXGvbzy71ufcjrmnuIqazpYlK0j5T/xc8JYlBFd0
Cus7NvvvZaJRzx4VPuLmqIQapeMQ18zk9Yb12xJJr+9hdR95HlcreGEQ1PsRNFI7ZFbV5pyf4Rx3
fWMQfMva6Hw0VJ+WZEQOkvWGpHslfxy/jVXtO00f57Id8rVuDd/FJRSMxMMcUCOSAJomEDys6pnz
3jGZRCZ+5oNjuvS0TH+sKbwS59lA+R/cXg+Pu09J1RY+/nQaK27P61jxj7clGcw2O4NYlMjH1TEF
74a6FLmQqwgzoYkNFSZdfPV2PJh0LkBxyfy0UZr6qhG027TivyC1lyQYikGRnSWkSo5jEf/t9c92
vy0C3Iq6MGYXX66U+cf6mktOak+FORlWARJ8iPvG2+XP0gHwUmqrkKDet+37vmp/PdqVo2NrAs7p
k3Zk7sXcILxAG/c1SOFoh6zamrb4Cpo/H8vzhk17KQ3lrVw81Hkb0cLnHXuQUgm6Mlb8AZ9xLL9o
huAIhqN5i992Z4/FXKZrOpSrpEGN0GobEB2RxhcCcbtVDxK6aFZr9bjCzUX//LZdRzttcPvglRJD
sVBZVmUqCuB/d7kZ/DdPgj0t6d9T83GbWIt/t8dasAG4KNz7qrlt7VFKHaLTAXzsSpqlJjUhvSzP
uZ+lrvutoEK05wmh0n1BjqGCCjb/OMwteksdm8Uz3jLGGhxPQX53QCpcC2tTOoj0RpoFMhON97Zi
7cneOC4t5FWeeCSFS/8XRNMbh115b705RX/l1f4kCvUyGwoyeTHYV571xCzbtBFzEcmYYy/yIutX
5IU+igzgb1YUq6Y89AJKpEF71LbdzZD4bwpUgXcGJDE0eErJHM3vFHNDFIFlebxoK/e/iwnQW308
MhM4VksfQhi3aeuun2i0wmUAUPlG0uTTJFHtCdo+Ij6m+f7H116daPRbWJD0TQ4rzAeTTYiQxL0h
gZU/39PfrpneB57yLo5AhJBASB0qYW+01FSkiNABnEmQGnXEpe86PuxVmSjWxoPolhYnBsbuJHtI
Sk3jz+coNkEqYH7141gaCxXiHMSOZb9+KAMbQu4zMVcTMRNoljHNzFHZ37moXEAAHq6v82k8S3XE
BOiKDi/zTQQogxB5eIyQwMC6kteiigshMZCNEHMUuoFq7y/8e6WA1xJxQni2WhBRPcJ7b+DcY3RM
UPWy5yAz4+R4Ma/9q3RGsipwGZhRb0BsUBtGiUwWJP+pGX8a41FtUM97hvWFZXvUCKl8qEi5c1S8
mTS26p8baVCaWkyoGUWhMMFRaxA+iK9umaLHJ65T8iOn34RwP8MROkD95dsdOGNjG9M8F39SE6Ji
Dsk0M+Wb8IPuiEgYOPWlj+oOAYdYkmOfhmuipzCqwVaG4hej03jjaQhiYLL53d/Z0QNmoN8Gv80b
I7e1T0PZaYzJre1PW6MC4oi+oLXLA4tMoooNyJr31v5rRKj/Zpe1iI/4NJ5N9E3b14y1mh60wYgE
BTXMemXK6E7g2VB7NUh4QSI4JxQT5P4WH/0S1KoIOW9aUp2HhFEX9yXhuqHhWjDfRBdzw9p0hjTE
Ho6q0nhN/NZATPvELGsSY16uuisGXdGlS8OVcR+z76evtq3Q1EUEViTx6w3toZatgIDeYehi1bD7
xo8INKAb3e9QZ+KOk8dvCZCTmOMD+nOgBc4d9fUmvHHIaBGfInHN/N7ti6GTOsXqOq4B+XlDKM4u
tonqXPMJuZD1+Auf08tA9TSEOKiAkatywi3PCfiibOTLXMZ2Al9uq6Y+0N1UjOciZHWUdccTb0wF
X2sIKrrUV90dfqhjFiVOisYdxfzPZ8wl9gybpjwmvbEvlr4h8ZUsCF3CmOM1MOEWU/3OGwHKAHqs
HzWKNOlSnDsIP6Gk24wXYL+dRDJjEz950ZI+rJYCwKQvYk/Uh473mkAA/e/zU4r5JMwE3t1ezZZn
kt1dV8hZOSpfMD63hg1d2bcOSVPe9rpYzdOXVrN/5BlbJ9r14qB5epZAfrGGArSCNBMdlKTnMeLi
sURDYpRli0hXVShou1pBwFOuuiMfeDzJB7n1PoC1ZMlnZoNkZTxh80kIJ2xtisWLT5IbpLUCMnUa
L+bLyGHQ5u1JadPFR9swKj12dy8tPJv16ZFsZwd+gG3bt/c4IbVZWnvo4t7ApV9Yl5fmSWJaC9e4
lK73CzH5qiJ8Kl4JFbvdCKpgvbGD/cKu0x86J3pAd+/QkJGEQqkrxRmagdSRcibjsT+VDu/0B7Ym
d7h2R2FObgMEUPP0NYhyF0iqpbLNadzG/GcgnGwtxCgEKKhewKT2boq/CRJhY9T5y+0j7sray3CR
ebgarnsjYWapZmAGsZNFefg6mKI8GGzDuRMQRsCgeabwCwGQBSdadLX1u4PLSnVzQLtaSvnsAbfD
P+dFX3OoGfmSegbVoA2vRI6s92Pd66EWq3yGj4yM/00VqF51I5Sb1iVN4UwiVYx4dILnk/e81mbE
Qd59EUwxAh48E0B42jIVzmcwJ0VImKxLkj8Frp/Y7WT2EOVlnMlQ2NxAdZN2AXMWpVWn8SbCl2L5
obj1cpGLz6OuUJEqmvjntBxWcFTTopU6ooNogFFfyxNaR0/YE3BhD7Z2BPoMMDne9FmrrqkDriDS
R7DyS7z6mWM6SbG+77m6Ptfbf6+eNVosoafzxjUK42An2rIQscag50zZTmKurd9KlO9T2bx/MUjb
BG2BpAh1Ak46zno2jbFazhT/Fi7i5T0ePTuQxsmDU43rCzITy9yN+Tq2Jc3Jq+CQyRIs87TqWDp6
LF/VA/hyWP3kiejmNICoMaoofy5LJkvabAY7La6fs8OG5QGhRlN0wN6uDkyzZUHBxZtaRoWZB1G5
7BevW1pLmJuLMy4QLELJMWTrSxHieAM8qXPjF4tlXGLFo6SXvneCV45p66KaJnazj+2AN1zYy5+t
+b8Gt1c46ffz0gBaZr+Iewvu/skvd6xH2GpkXaBtaESGGv5b1PEChrY1BGd4jUxHrMVnkhm6BNgB
Chyu0Eeb46mD/NSlCwrumcDupV5zEyWw9WHbUGQ50nVu56ctDIlTIeJ0/muvP/tGwjtqZ4QaKjid
cYi4KhQX8+AChuftZBGzfcEQjoEZidS503qHw78ORzAvZaK6kwmIOTpl5VLP0gydmntSj6u+9DAA
08WS6/SF2Q86ydp1gwLGqA/xNOqPh2wKj3IA1X0wDx9v0Vtf/2aXShbMHABjZ4FIeMmd4D/lskIO
rxdSllZFeq8oDns2elV6EBIsYqY+zTLCsnNESn/so5DTQt6S6LDIdsiKn2euQIJfatX+kcSaySgM
nNXoKe6po19rA9/Lr453yqUvvsQSL07aYw/YC/o8oLCfVPnABtZjvmbT08rzUuR7w2MaX5jDGiWO
uhljgaw1nE6C3/M7f8mP+Ex8KlgVZ3qjjtmhTJTFxOjELSuh9kFmgu3ec78jQVNVH9rFJIJc5neL
FUtpZQ/qXliRiEKcaWMdOVVyJv76EH5zHNBO7Nx8L/fMlf9zSds9X1vtdUSQgcwcFxxMqIUe2Tbl
fiLr7CELSFDCr8c/nIVtQR/9O1WOsAK2nkEAuMisHXY1bG9Ay/KwR+StzVaBJdJK2RkavUrzSTLw
OyALZ9NfJAqqwl9vQEoBkUwB/belD3wowYLmrnUL5YRDtm9dYYYyCYQOTbOk4FKraf5NbzvNOQtY
Fvg+DevXU5jcAtmICYiK/klY482+f2Mr8EHUB/jjQPSmyEJxNDF1w+WFhfG3Mz7my/KgB/v2U/+T
KsVm8JaEwHQasCCvs+PvlziEGnQ77+rSQryDNvruq4zYhW6g5We+rDWLjHE8egTC4ep3gzzRYegz
Mb0MsZ23yvMrYDS9CRwJOs2tz3y1ifcvYzZrB2hDKHBkB6a+UYgh/slexsgYuBt3fEHlOdGo9xaT
AFfX0+TGe8pWKne8U2jPKoKvTu1pMyw1NIS+P3xTgVjs+5Rs5W8egNhbRs8kThcpeA/GyfIP2x2H
lz1BgG4LmTCEi30LI7mhMJmO/+9PK1d0/hINQ6TGiqQn3/VolNXn4YD4B10I6I9Rb8OKxoeP9c7r
gAJfLp9d/p4QWk7eEzZqXruiuoC52sBOB1Gj706/V+ML7yUg9DZVGLSvEYO5vtrPWnil2/XxBRZY
FitdZIhzAzMeR8UKRoITSQ+W7Jisrhrd1V4KThzK/Ycg1DVMSqymY09Q8CCd+PrOzLv1u85x7V5a
plng4zBvFAjguK1X7b999tSkUTvGLmRTPcTe6z/MU5INt3fOYHtL/H23lQ5z58QlMnYmKxHxPao2
kzFdnWtg+e+xqhRE+HxPKdImf4YVAuKpSLRajMBAvsFVsPlnc969ffHFB7BBaRMcXMwWyBS+63J1
4K1oKoVmsh+24PPocMvlqBlXhy10MLOaH2WR3iQfm5NQv1ELRymxJmwF4tGxjBtF5wihNG79GqgK
wqVoqqNF5c/uJDGqHyj1wqNF1PhtEKB+QCoMbaW+lbwTedx69Qg3YCxSjf7T4D/lX7fbhPSqsSae
EhDIayo7Gm7arNHcpOgEuFGNmEPKbtly/nptMU8XtpPyYAWtC7FgZoW6rcWBWW7nHop1jImUeTmm
/DL3RcL4bFk5QdG+GeUXab9d9T9SOyHFRFU3MaQ6bHQT164h3UiEen91aA7KdWYFfAgRGch9MmyI
Fho6KJu9eQ/+RIsrTCdyEuWf8xlOMSQTdogCxIeflqioB1M5S/L4qdTCPIvfpfzJbQNZX1P2v2MZ
wS5vgjs6Kya4HndfodyKr6J6H0iTuPHobe5BxPPZBW/DlisfSbMxPNQ8bqoNdH8zrg49NWRqhyG+
z/O8f0R06EQAujTOQQ4wwSNzZxA9IEUfkSJEDTj3pOUc2Boqm/x/YnTnaFjmWXX5rnEF5iSUDBAY
PNKGEv1Pr5nzyKp04eaSNbamsn6Vr82Jw79cInpAAGhU2F0AXN09lojjctXZTHQ6FVJUV4iX1ua9
Iz6zum3h62bAd4AOf+KbkSelH7s8Sym4EhOKgUWkpvpv9Ym61ClLG+QMPw9krsC1k3FJCaHp2/QL
4pw+YP0lfgCfxcEcBlsnycMOAXVEWRdZVScEI+7Mv5eJhWpGv6gZXzB1+stkQPqCynW1zrX64bFP
U0LxM8mU8ChoiBo49a2jeBC1qHb/4FhMXSkLk9wnyyXQIPOWEwdPe/FtN9EEA6oq4QMJfikuMws5
JrFyzdYyzh17FWKFjCNef6UVPdqAWn31LvPi7MJRoIXfJTJ3XHIol+untHkLnyZZ4F+Z1EAwNWTq
+TVq01FcVnNZaKnSxg3XGYVjBWviep4DK9vZ438FjX4/YcIOktSA1fCuhAjK3RNnD1uDtv3ttUs/
ud0PWuCxc7LhNUapdCK2uF0j6UrIfpXMRGt8yhpF5rAqwG9QCFJ2vFopGDpWQkX6wLX1rnHFhTEe
5rXfxrcDZqOcU4mCeI2ESqhZNbMOVw6BM7B6hSNuALQ6vYx9nMyOypQbuu85lGSJH+EtBsvJg7cv
1SNJSU1FCPlspGAujcUmzCJwA3fU33TUJ3NbGfrjzUap9L6bDaWQps5zfZxcyCokcMJr3bEMqSfp
1Ne07tPqUdAlLwUrLVd0DUYR1qQqOCVmWNVuWF1aXpvyrMOI1+3Vqnd016pHVP9KP6EqtK/6VIA/
CK/V0TfNr/qbDHM9ClUE9sqwVTZeVV+HbL6a7SOFrL6B3ZKvOWCLZznPXbb1U/gVTMOa7/02PQm2
9yKqNG8aQUrTa3SnN+fFUrRPwq743/1wWkVZ1dMCukB4N0Gwm+INAFms6EZ6Sgsg2mwx+qhsk9gO
5321FkBZgEXdMLlXhnqJKwRgY2cpjMT6ieqMG5bpEUjNBI31G40MmN5twu5uu4ktZLZ/NKsZARaz
WyrQiiPTPW/vILZzyaDa8AEWiC1xiSXLqww86Kn2YrxLrZ1hbgs2u723UMP7NyyQWAyoQX/KAs3m
zkAG5H37AI6S/rYgLPhPjpLfgi2Xj55avBXy+sCi7M4Qd4IYBlMxiyWy0xXB8GE2NIUKggHY3HGj
ZTbsMpchKN058+2yuSKxVqHl0qSB+MdFf9/T87j8LF+P/tI6daby9FEmObCZ772evweL49ukLdxo
+FTjT4SZFyNIJbxgCHtHKBr6fRtaWfFLsS4nyEuBHXtoiZNpawlDE4n15m/ojU0LYFSaxPmQaVhg
q+id29JMwe9l3zr3bhzSQZjqLB2NK/tquKH/JyozPwnccoOK+tmtYqXv/o+puBMRXqD2QEdl1k5Y
XFUapFkQjrEvIX7Mvop5rV5Tx8LShqoCQpLLt1w92cVD7d8IbH+tORPMZweO968kpwo+AifYIEsD
b64rrQ1ta/e57BxxtdpxVl2uE3Zg7n20kLPvfjWb24qWbboFQVYs46FckPKIxDeWy6TykjZFsCJL
P0SuGWjN84S/aYi8ZVR1681RrDvrSEhLQL5790LdgMfISezqkCQDQ6Epf1uMs0wNwJPW/rw5B5hq
DmbgwRq/ujowXH8gbbThX9n8sE+DUyXpAhkYaOp9nCv+7QHdnrtvF9PP+xhOGaHbSo6EUv2MT1AX
eRyRcqHvTuWvKcgBgOk0xL1R5OVSdCv4Mkq1rTC7zl6qpRjVuyNBR01zpa3kEMci3YsHVekFbjOB
EYy+3qiOb7IvwZda4NQg0fC2gFXpV/ZGyl8gd9wljh6L13DC5PL107mxcWCIjK3nbGodOJd/nWG3
dLoeCqN6b48CY6GQ0G8ndM5/Vrt8jEqW+gK3PmxT+0J5nZEmMZHu+XLWdanFt2YKWEMZ51X32i7L
BLoaJUTXU7Syh7JH2LR2N+e0u4D6MY+Z9hRHO3IVzj4E1LT9MKq3NEWHrubhbZny/Zxyp46OhvXv
WpdVgwrjJ61VUso+YKDEhjSPI2yevjjRPo3HRLTsXdtZLL1r0uCNGSSbybsTCCrMXC/FrWFIEjr2
mYPPllT2PGJ9Jn/gSLZ7TZsW0WL/Jgk/SK161b9kL5bEas9YD+UwAgEjzx3BHsWOBf6VtqpzDWy1
qADAY2iioBTHV3QzVpDnsI5W9DqH4T0SsxhKjVJNVjfjQc7cXf4kS+95yP6T7+/5NecKmRFKZx2e
Q+6hHDzvcW18fOWaBuFJo+563m3AxXFEwZc4WXozFl+8jIAZgAf5xLeUMHhazlyXS0YDDcbEu6ju
OWGTQ/BeImuQCVzR5swWYkVAdqzh39S3NAyAq7Q0Ac+apfFhNpq5prXmi67TeegnpdqTdc6gkFRi
CGHpRHGqUpdX9uz+6wN3pmltQfZDUTi3+ZyhrvGGifvDopmnMjQDsDyxs7DtloRmbYGdvXNng1X0
HIc2wjSFQSKL2TZmJgCLzkJOrqZO9EQOrFGSyHlRYXtPdM+UCXKmVLqiISa32eXc3T+f9XhB9mDg
jDMwfmbF3OG3+wekTzb4r8M11nyG9OA6QDbvkxpi0I20uh4zFBegbWyZSAuDrFDHKyV8Yzq+iMlu
X6Of6GRO9l01bn+p5JYxBkzzLvE8or+admoiqrWhxV5mKfMPPLPt+gsMgL/Xr8u171+m2ccXWfnN
ZiK/IEuzIyeGgxoxxUjurBgOwkMy5eAzP4d5fGupXweL60o382YYwfoVUqKzht550+/PJbooC3kw
N+BrWyt/OnaROJd2ffiMkuCNhKfaBC8VFiDjUI6lFnhiv4WdRQt1dyT8pjb8EJXPd4nM3AyBifZZ
tUKqcL4vBk5xWWEspyFCCwMM6BjD1Iq4Q6LwqqyJzdnHGyOdojIHrUWCnHm6P+nwQ3Jy9goFXxlX
CwSNyPrPzrnlWP2OLkpIOYBSBeYRBzdXGCRi1r084kn9QjoKudPktXLYC9wD8uZSwnargrOeS+S/
Qh2F5JqWFwReZ94K275huivNGyJpk07HBQAbj50WJvVtlzo3T73tnVE0ZZ40wsL5TpjCK/e467og
sorVUOWM6F/sob6ABfjaxmyQ10v2pfr45yRvuIVKqj/NXZvyaVqyqxA9ehpOJBFzF2YlO32pO+yk
FKDcjjxPDkZZHuEPLhVBAzVVn2oSwHlFtU7YIz8KtxiHo7AFwdqqXAibI4fuSfK4cvjSU8LnEGaK
TGYaO2bYSyBmAGTu0JojkHztuROurtVflhWTdEIu8KH8tAd65xPkXE6GlyuIQEhDMbqK0VUMpwGl
7fAnHB7U5GxwqRBzfNg7ki7nxfWqDNBzmroteBM60VfcqvrezkovZLHp9CyapP0qoRKz9nV3zC/M
qOpf8qzuPVXyiQof28B6om46EKGbmtQiY3K0Cfu/nb8m1ZVFXcCpMe8QzJVANamxZGf5g8NF9ZID
xHgQqmeaOD835gXosCISnm7aSscu6dkbP+0iAnLVKkKBgiieuu5/+l7cKCbMWo5sWLxgGK1RRrow
KmC588eamZQ41xehqTf7bHm+4iOGYLqr5Ll3Mv1ZIhdsEgGizJWWtmIU6O4862m33QZx0KZsDUb5
dpMKceZmg8hh3bu9CwmDIhZA/C9yb19Bcwdu7q6+ZBc03PZZtO8b15Vt/T9H9zXXjczBzHoBO2am
zvRbrPAc5o4gkorN9Aek6DODjMu3MNmqEjgwsihP8KPSqhvqI1XuM3QBBJ/FdPse6gFKrzPUoZqn
CzByhLtwGS2OxPzPVgm2rFA6tZdBfHhepc0Vp7Fhjxa+b2CC7+DTgPzVxp8HiUTp7F8eFyHkKQJt
I7ozR7UvkSXHVeXekEitlXrDQOwJLW0tKsE1/1RJBILJC2dMxp25tplt2tSKyxbQp0u1WVZmDPyZ
eK1mv0oP48zgZUmIiAbPCCX2tMTkpLYAx/KQ/Q/mugy0jQz3Mdj3FHjTk6KTFCnlmyO6RBjfxw1Z
zu0ZEJ/XyCJW9np6L7IDAMWSUfz35rCqlTZ8tnfE/7vrLFhhKMhH/J8IDZWhoKd5Q5UheHMH28jQ
DOlSYwMLdZ9S4uHX/aZyqPiynoDIBFw63Ip3Z2kD07ZrnAudqv2pyaz02L1Rr7qfmonUEs1+4eqw
R8/M15Sjvcj20/vqwFGQvVXQ4yhyV1iU9dSMNDW8rqwWco7M+YLcGgPglmOxim4en9Kf4lpRqlXf
tpO/FYt4HaXRMcsxPLNuu3S8ndoYPemSePOBnHRhXUm94/ELlJaAHVhjN2YmGGik7CGX6KZgyfKd
6bRT8hf4uQULs0hg4nuuecUw5JK7F9yBKOGPtNMLKSMRuCleXvcE4ctg9WQuJD1Qr2waLRjEgCEx
YhL7jj3U3X8nBA8Z2eOUSaPNN8sVv8Azn/YnCe4qEmvdR4W3axMtYLRbkIBCxA9txpAAuVPPdKeR
fwMY3cPj4XBlWN+38gP3+Q5a1stt6Tqa+3HBkWbiRur6s2AxJLV9UVJvpO78Wgux2cgaPBw2kMHx
ZShP+NM6LXwFA9Aij8DmFbfKOx3b1zVim7XLxpIZ8cO48z5JqVYe6VElEosSxuXD+EISbCtO8qsD
R3D8HkXRUkthJkmus4s/LcHhgQAc7aZJp/6iT2/dlQjTgDQpxXphefH7kINPNlmo9gfdBQolQ+5Y
cdzARNe/Qtc2AY/umXQIPzJnzxTx4KU0EdyDJKOyrM6lnomRWuAN2Y7aQZaEuhPHd5bwq/hf3mn9
TBGXUyIIxzIKJmF7y9YH6FczrinWdae1F5Pkedz262B0XCbakMu5zgE/tzH727GVHEDXRJf4rJsU
3XNfXV/PIQtyPjbMUIP/EcUiTI38XAc0rxwwbrJ75IK6b6THlkODuTMO5hBjtReCgHi6T/nwSp6g
fYhTvu5ZLZqMKuRtA2T3b7JQx4HIHMDJBWGMl5Cj91uJ1107Jf8EXF67XcpoZP52nzYbYZBYkHuH
zD75v4sx8NpyNtVVg60CE2JA6K1WebWu6IhA1dLBpNMpeIKbPQYjQ6cNI3G4s0D3rs8vRWaA0J2I
kZIrAh0pkpuIhvC41T6gLv66f4vKefmJtZGZT8917ntSlCENlypHhwSOEwa+/cAj/CbTC7eAoZ04
7cVLZbP0SIbNiaZ3SUMoWWvKwJ0kmiGadJ3kcJCGdTSe9uELcXezSgLyNQqYj6Wyfi2Sb24Le9bF
Ui8Av4ny3SD/9ENFjZpGrJTGJ0TgbZFyW7GDIcqeORyvpF7e1VLui9rpDHXcpPlE7waipupY4MNu
M9X6UL5iLxEKqpeXQcLvo14zCBtl0/FnF55YTnPhM0c+AFNGvv1oBZ2Zg7zV6f3kdiaIfot7yU/Q
IXrvF+njVEhxQcXGjUFAIz16Trq6qmgvZjhE53b406Hnyl/quT9/QpsGXtYvxebiHHUpvrfsmseL
shKuNsYV6u/avg00AH0EL6HwrEjTA3XSd/dSLqAEannCytLnKh9sN7BULrNhxSxopx5wtPfPjhSb
YwHaSm4kKJgvI4TEA18qC6SOn+i8PCB2tJ9z6+9ZqZsFIR7Jknc6N1JWrVYo3yPOETGIZ4at6Zoj
U7l4yJpX+aOlMbxcvFWj0y31CcrTq5n+gGqskIzI+aLIeF7FRhFTVY2LKjbEJOGrhxurE8dwQ8Cf
Fmf9ULgcrB8S489Iziv6pb+BYa0vESteg7zqVYujIiMqd3UThfApEWtfeJMITKLhpdFIYeqAvn8P
tq+5ohIXYTXJQXwclq0IjlIpGnyKbFYm63qg4XsvyZxnac0bseZu7oBhpL3swInYAhJfYAJSG8nv
sEHbPmicjvboaoXy2DufZMNRPLUKR3fFTzSSYlBRs2nvluLP3dAGJScMwhiRYuK1Aa50g99ply75
KATU3MLYPFVVTXHovW6hlQwOUF8LV3Hi1cK6lXI5oL2TWpzlpnPzKGxPJN9m3SYYTQa89vnwq3E9
VHHyvJEKqQIVgYsL7iYVj1PPfP0o6A9pC1nA7XsrsmoE93XAMQgjoLc1WXhp5u+UENh/ig15WDk8
0aS0CrOf4vWfVg6n6wNrfOYX7E9+zenRPPgL677H3SQEYNRZWpBzY5Uny4b7Ppnm1suullVXgmC2
sjsDQZFweg6spBbL9FCbVgGJNphjxtgCmrvhw2jgIg4Yk9Yl9/8mqVHyxDnKLMioR/fcWuusbuu4
LHSAWTEdc7dxSimEwjet84Zwq1uD4OIvbdRm3Vo5P4qXIFVvKNtBB+UkyqAr3y4oCZSQ2Dt/ZSXA
axuvbs5tZj0O70duPHNvHSkMGjHnlDP15XjgguHymLvU6r2GGFaUxDEDzjmBhMn8FzMgMKvxFWmS
zmk61qo1BWCwsa0IcTIkaFUJa/hNn9u4liaBjE7gRrkDRHc8tq/w4dLnY6WoJrQDy/FMBu6/9quF
+Lp9DDv6E5kN+Tw4V7Z2dMriWye4OV/PbwM8HUhOwCuv/ValhEKwdcYY8uepDoqEYt22dSp4qfk4
NacnHBj93Lqa7+/LXFEXmT3NUyp6p50jB37hpMuFzXjcmY2X4GHY2rtZbWZN73HuyNr+xbfNKIGs
njVfegJxrM+S3XfS+9ZQxNkkF6G02g81CTLx/ZZtdBj9k/jv8Ps6a1F8pl4WbPF4Kxb4dO9M+aD6
6VY7x6kz06cUfCKptslNpesnf7h8cEhE41tIO/522COLT2EkybTcv/vRQ/N+Vap6pzUqZR12CF7Y
25G41YdWvdMXuH3Y4JsUYpCC+/7DP7utCRS6DSLr30jvM5V+NivZNNWmynNgHJsTfoR2svdKnPHi
/4X4u4+L/z+BEtncm8fxCiYSuf7xFHxDb/Zy4hNZAsYlnnWl33ndYyZZguYY+VsOYAmKGld/ZAuL
viWJTwqhZ/9ReSKwAVhtiYuGMkdw7YljgVrZrLp9BaabeRfp3exnSmnxIzEFbZxG9mngYpUHpkD3
DGgm3ZJmFHVA+hHJnGZ8CibW4kLAosSwAxoSxW23e1Slghh9rM/T616UreE2IvBJXUGG0XbviFce
lAlcFylCcfi2wsirNxYmLCb7tBNnrj/bSBY155HeCb+prAwK48u1bnQuqHOMbxeYWIfGogl4CXx+
Zz06Ybqum0ZHgnyD9A1f2iuKDWhk6Ttwm/YfDQZyHj+a2uEYV7SaWbg53Q+pGQsDUhzPq5c0Eo9g
a3Db7LJAjVPfJoTIs9yTNu6JrVPF1+Kjbr8xtVWbFxamaykRd+ynaTbxTnnbD9d1gcBdujvjEV0m
Or4NrlaGGWR5O8ZEHJOvADRyTg9XPBbj/RuY5YlhNUOgP3U8tOAW9xWWkB/Ja+5aSv4tvd3ywSY/
Xhq8zrktoHbQFVOFlBUcvUt3xEIATPpBviBCUO3nWk6aSSXsZ+W8lErQOnaCsqAwSoIUkBkrXE6v
d7O3tVRHxG3TBH8bYx4Q+stPGM5CNxvOh27ZMpfQljzeKpFRkPWY6L9ShsygMxR9roN2kSR2Oc9n
xu3DK2iiib4X/qsVpg/IwekNU5IkARRjUxTJLQUzFIXLGptOZM7P+89piHgQsaD74nBWfQELJ3OD
t6998/numE3PpQ2EuK92yJhs4VS3wgHgzVDHdw62bl3qUFraACND6ycAz/mUy+Gx0f+jPS3YqdNS
LfxOBuyoVCwVuq5pW9nTOk1r2ZmsAhJDDBlyWanXfMbT11mgefT/D2K1r+T5ASZbsAowd4Nr9c+U
s8y6vKFGGeblFLnrTlHX/BO6/HusWZu9RQnqVVFqpK47A0wL0jW1wLXHPqbMMJlP2hyCAmIRLunm
FbgcXMI65V2tBuL/h/nXwNRSQTN4hhZcX+yyyQpLrGhcpXrXxOAgdU06Tcd3OyXn+ci77R0ghhpx
32VAQgGR2jPlmDVEsijcBOrKE56sX6OkMwZQ1siNA89H/kEj+moz0mbia+SfEXLjWMNHZpYpfNXQ
2skAZvpRyljAxJ/2E5A9Xb+gf2QRDVQZbbMyGiCxyuGrO7w0s/xKGqkfBMiIKocxDISK4W4uYRe5
hS3dJxOX+eZct5Akjts7M6y9pVf7q7vGi8abk1hLD/kKdYsMt9Namy5S6uhk7t7BffTWUQdWWiAu
gTtuelX7BOhVPCUlMcw04ffrRhypaHdT0yk55quEM3QCb9bDosjLAN6AK8XMmuMInfOi3QEZsKmN
2IOL0IG/XBOTyfu3ume1E/7pJz6dfcgRuaARqkGw1C/EbIA3594BQpqhdrjlND/I5ylYvuMhDAXj
aAvGL9ZJ7qCRp4+aR2y2e3DBba9CpdIy5EEDZ4/yhtb96bGDzLusYiTHSIuMCz2YDlH+v9DDgfMV
s8G52rhSbNjJI9yewBgLGu/HU0R/JjdLKGaLTHo/mlsAvm8VjQwyB3t07vYzjZRAIVG2PGnYGvVH
lmBalQv4Y8Wb2zk3JBSxyR83ORY77bzp8GOeo5WUX0nQrTMv8vXAAWhYAzW2EJ61HRCm+sdNd74/
VfngXmKmVBSmgDbkl4WXGjx818bHkhbLLdSsJ3Y6su4S+znyiIpFL9BYlJ5GVoFAocqoe/XoJL8u
iL9Kl26bRPqrM8ySfFB+NkBScom7AjSZvThxoiJA5Qh9v55ijdDA+gScPJxik2V+cUMJ5bo7ClpT
B7aqjlRTjhUiAZtF43Fhe86UERjvPwgfjmYZWVTnTt7Fl5px6Sf+lenIhLq4YHBOmR0Tt1d1ylv+
Auuj145KCzegCYUTqZI9IiV/frTX3S4gclLxTUhupW1f2qVHUaUBjZvSZ/wPQsYthNBqWiquOrrT
N+cXVAYeiLRXHlU0NHv1ixPBdg79deDxYvW+MApi9a0b6BNYqA+uDZEgThV3YUudHFsa55bEjcAR
56qZOloNXrPktWe/UwRzCEjNJWNq1+SMTv2CUOHRC0j/eutz9mzzOFInjo4dVHS4iq1z8qK2bO8Z
vUuusyRBfaxjaA7NvgwS+kq3/GRdTmjBR90G4pz8tSAHOZkPVoje0nf9iNnSdriMcprV4BDhGp5Z
c8Cow03WMP20OT5CccIJepoC51kSTCuTH5zUtiduCq8usdRYqbRRkmSbDgAc8yQbvMp0oXHhWOza
Eg5fdac8G2jPHW6XZQ8jEohbRm0PxTbxfxS4NBIwnaSVkgfAmA2LVSsyxWbs0BXH0kvrw+TZ+zKs
k1R+wtm9fAmtbJnUAiO1OXSByyK33yJowcuuvtFD+3UUzW4Pf4DfSVEB5hXurFX0qk2yY95Z/Ok6
mk+yF/mNrEp+nqYU5iqW3EAkKzngcpZBTJJHZ0qMcolHEQg9wQ1XU/bafuIDiXIY0bHeJspbIOgE
1GFWCVi6vBrRwzG5CKNoAyR3bijTUsMZv2YaJPPppALeie87MZRPOPgIyUoLZKAtsb/wkHzcEYfS
A9Lt5ck7YRHR126gEf6lfmm2hYrH+H+Efb9vMtscDZf6vz6IYftxQMFJOVc9rE15jOhJTFjI9d1F
XBxY4VbzhoBWb9DC2Yobib+4BaTCDExWdIc44NciLVzDWhV1av/QBxAK0OEOl9a6YdmCTEcv30H9
Uy+ixC3kXyN/nH1Nh6xqZ/3vck8ggZ1VUZPPY91nCwHofYxl1V0j6CcoTaUIQgzKRJoSdbf7KGuA
0mi8YQ3qNYfOKXjC8m+kyLjAa5G06Z3kZJ7f8ajtejbKbzke+ldjGqnMRsaUz2YCzdwvEWlVHdpr
j/DDxGb6ROjf8Qsbu9E0RD25RwgTYPvNT7ghQV6vCuMduwWjw1SZC40SMLrNP6RqA6eoUvypeTpb
PGhJD/l3Eg3TxiQ2L30MRF7Ky6gbr+8THUFa2EaW1AWJEYsdK+kFb2YQcHOSGb2X9Fgla0jGTltb
5MqlBXEq0kdRgZxINp5Mh6Otz8hWBCjdf4tJf9SfgomTDMZ6rrIVSaSE+35BBgvJ9FjZaRFVKKKa
9FWPJs1pjU4SLvHljTwZbdJ170S7PdV7xgw/LzgoX+muLaF8yYxND45QbTpx1x6ivHS7dg+clFSa
E9phRILjDCjJEmuUPN6LIrxQAiTS5Eh6cjWD3w8erOLDs6G6MtsWgcXGLBI4yAr4LI7c0zjsx08F
WGSYP5KdMreBdnHPjZTDpRUGiJ+OgNp2t6OvTNjm9/uWJIQzSyGmXrksf0l0K8fkTA+RXV6OiJFg
OVVpLtzKXHsgW4Y+ZO7cMAoz821d6LPVuB+HCCAnUsMAqOiwQi+ceU7usTD62tzvCQx6LMC3pRu4
1DVqjil8Pv+JX9iUi4fHYwwxRXjkdiinVYzLU5EM03+tJf/THBDlQYvd9dEOHtSZOBIvn4qE8q7z
037E+Sin+7ltHNCSi4kZ+iBN6s3DyyRcJFAjrgJ3FD6WUFQGVPCMiNNI0DTP4wGGD2SNTy8stqFR
RF9eIX+FT1BTquhWZ2tnSokseg8o6t6hlmyKclSpWyFFb5javKBG9hBrSsIcqz0SV3LL6KBMXFa5
Q2DJf08c2tSJXEEjawRS0Kph61C5rhONYuNh+14bF9uE3ilJ0bPw9ofo9j7FQxJgH8VM5w+F7Sh2
Cn4VUjj8Q0P8pmgi09F6FZKMelTnMlmQ2cWTvuSnzj/lsjUYYM9cxjZlgKySPbO9pmcdAV8AzmP7
EMoLsITgNyopo8ljLy1Rk9YfBfsEwk0QnJ2XzTcbv1GFnlA1pW53pBXzlxc25Ud6lf2bCcLkIztf
1k5Wz0xFv353069ZtGEqb6EMuuD7a9LqlvCtwB99/7O1WZIUgyN/8FbhGh8hN+dmeH/lv5/gh7Zv
GpdoPZx6FTYCHrbdGgDCIYe3CzltPf1OZRzV45PgD1YG+Vf0sEafV1OO2e4xkDLQrD8n4bRYK9Ne
pT+3crfO4yu2fSx/HtfcBPsFXVHgPng3XVkg5f3gX48oF60rdAcSQBZe+Gp5pL7w2KQYDwoNdsTI
9mSDj4ZVkJJ3w59KUoE04NlVDEmICwHFjsI/JUiiQJij9xSFfmIloYfrZKqXK1l4spKoL76dyIFM
1LqN1TpmwySkk5iZJB1CHB6u9JWiobckjpvDKRs5m/OulmgJyjvHAZB7B4LwWkWIFEf49Yc/Juab
U4ExXTlipvLs0iMBxdVFjk9133w59ERG1Irj4oqGnQNOwTOX8r0wP5XN1FzwTC7K6xl8vU17zlOQ
GPdSYIPiSSbucSrSRCSUJa6d22/Wxpj4BpviitxSO+26A7OI6m0mCmN2tKQfrPDdlXnEJzkGBRw+
siKEwYfHLSsaZXkBdZj2Q9S3TYTfIBbXCaycKQCJsSrJ3hZsHx8HHEVyfeQZxO8wIak3pB4YohQO
dL1FPIoHDrb7unip5XFr3cs62CgZeNBOan8sVGeOYvSTD8tFeNjURkJVmE2CuCoHcYPf0OwcnEyd
HRba2McCJUpbMxJpgsbgGCu1qsWvMtyuT8Pf6DOZ9pOkl+ER+fce1m8oSSZ4Av1YLjWK36X+6Gyi
nJRPzfCrXAqU0PHQWa5jjTxgy3U+kYRudOiZcSQZx6H1NuzzT8r3wKnSO2anx0FguLbq5KiB6eAF
ev1ZkJfPPFRwJmfsPwFJPbW7j8qzOzSHt2mFxMtoJvdJzAj+Bki4A6giws85lJB4cfEfzShvYkDH
0Mi29IfQAEUijrz2Y+sDxVMUOkSruOaPk5oDvq8VyI3gJz1vBWraKYBA+VU4bYVBcBqxHBRrOply
Wf76ItWf0oeqIzw4++etWd7NEdQ4Pab8+19Xa4iE3mzOh94Mhx3dReHn2Ljz48is9w3yQItIZFia
1pEp5+VL1SYVzs1TVOss//+Yq5Mpy+NXvdzpcrbZUQf5XEJHLl3T3cPrXAmeMEvbIVxwGzFspO+S
ztEgqEbIxsHo+PNPu5yv1FKRV3VtG4wN/ddgolNR00FptDwPWtWo4ThszYYyeJ/F99BhRChZFrPP
PSZwGeoOIkdCGfcGjNaJSyu9G3Z2Rq3pzNziCa54LIiiTjpwZT7p9cGP8+QYUXD9XK4DGaRjb1I8
4gdkWDt7xaf4mEA6qc6KY6Pp9wUliZJM1F7LeNgi1ifwPrW6KqzLjOMuN2fld2BI6qnDP3trOrlE
gP3RAyPOh4kK//coCknt0H07YuP725X3BbuBFIdBr2iJPM7ZfOom8cqtabNz6cA+tU2ia8XtHicS
fQKKAoXA2mcTwGeOLRHTX3ACkujFsrrt+Q3Xh5XkrKnrXiFoxWmUYtsHYQ0cO+ElW4lZGrvyqvX/
tIPLHHx7VbTSit6kjK/+qROEcIwUIH4x620j99SzFYa1NsKwvGciZCihN9uSr7dpNByboTcNS6zH
sdH2fQRhSqglEm+BFpq3mqeE9h1+scUF5hYMXOjxZbSe60JbxD4ZFuqgTWEk0/sDILcf2MiPbt1b
VYIqvaKmEZvVwQRe/Zq/ryIj2gkgZyiFVPQiwa6eBWKUlfo72sAIqFXYFcWfhZ2Tlu3JNaccnjng
zNQStGP/4Q8rA+ZTuvLxGIvEUDWUyAbcwZ2A9+eVyuVvGxI9SOFOu7J5hWyaw3XG7DYkcnJ4GabQ
C3WGVtmmwj613TCI0BGJaTbe+7oeix4E6ofdNgBISX7l3FjQHDE9U8vx/14uuER68LAPeLo25bkV
xJDmXEyXVZ6njqOvU6d1PI4qjc8t7Bk6KqWYFJW4AFn/dAPkHClfGLi48XOPYpM7tnJBrgkkogeG
WvCgj5tL6f7n+jaFgtlVvsgZ7MGm7pC+dmrkET4W2k9w/ChaBcYHnNjVmS/ewRMCMw8WT1oIpbXk
2eJcS8rHwk+oFsVgYuzjk3cnbsAYCV8497zPirCM7TpnS2eyyTVf962aowuHSVjPhiURM0sXUPoN
+y8nPmtmj3v0FEqC03GSXHE3S/sthyB+Xzs71BC/mQ9DDbzw/hp125hcotSUh0tGTLnpFbDHwABE
14hGXzYt1ERdpaxuj+TSm84T+1eQMIiCqHYd6WhIBg5tnGfFI7j4wflbvoUBux7GJckj5WNno3ef
hpkDFf2T8bV8yvKkeYmLQP740fszxG/taAbK3/ynImqH530+w/0KzaSHkzCe+ed0+Mlu7CAG+14q
arlfFyGYPUfGgml1lsnIR0OS0k44sGlfLVo4DX4GSYweYY/kiBeE6A4WMYxRg7c45JT6QoY5xl8A
2DK1g+v8WGdCTEN2qr8P03gPzjzr85RFbusEdqMkJfJqi+X910Rg9R+aqPh0u2iEYQGTGjC3zqyW
CgP1aV1tHOxMUKQFTFc8hX80ja6yeslgWNVR7LOO/62cwA/bEbeI3cWCpqOCVmvPs16AvqxB9JrT
p3dOvwlR0ZejVVucfLq8i7bMkwvo94JRe9dNdN2hbDt2eH5kMe3kk9stBY7MwpGpR+VXkx3IgU3/
+MME06PlEU6kMnku4GBvshhEQk0mX4jAckGEYOIOF0cADcVEAvDIpq0x5qCa0Q8GrK+GX1gNRJMv
ecWkrtD5RKKgZdvCtudg32wdlXxcgpN308TynYr8/hJz5w/6wye9WXJENu5koFZEJTtr8RtdK62A
9wu3RgnXSS33gUqffWgrkDom0lhZ/FP8NetIz6qDI+1XQV7VXc4mGqMEg4kbeq1ok0Wi+Fa6Kjtl
izsMcfEofkod5j35UJVx4y9bEFSQpKKoHk+7TcazYfhVGvA650NmV6pZ++NWQNX9KDknncb/yatZ
dHk9urKdixHvZAFpWXEdsba754S10iP38UlD/jsOinQlkF/BgIzl/CVApoItkjf6I4UcmodizkPs
NT9BsZf12/pB4jKT8upYCWxfmtb2FbEGGl3ysMWitlNCjPulp3N1pItTRu1FbfdQ8VUkM5rwHZLy
xVPCOCexnCfkSyRv4wbfTsYuaCMzEBwGJ+6FtzpS0XvgeEnG9UzTRng5p8w5lsmULdKXzV2c+frY
lsJKSiKjsAN2jijm/bN0dBqcJsryxvy1JpAqr31FtYEHJ6hYCWnE9sow3Q2XWTTsjbaIB0nuLzPm
W+p5sUsUvtC1fpNe+FTOsX5PchnBO+joem9YtrcqkcD+zgw7ITwF3U9EpdMc70uMz8K56Wzci4Bg
CkRn5nAzr6LwFJn3AIJAI5SilkJ3IGSNrzvsItgT65ooTuqffpQloTZizW0FfPU8ri/f/oM3zGRj
D5Sv61YpyHtWZV3hNWXi3afcjaLmr2W8Ox6HMt8YHUfRcABN+mRId7rlcpYSGe0Bc1IZ5S2octfH
WMw3Tcw+iQRIFNu7061Epqd91VSRExg1TqL8ca561SU21a97/foSQdXMjdYrsk8tWKNoSDLMAkLr
JCZHLa4XK1sgqyhPg+DAweyC0i6shlD4BOD84/C7OpRV2yt84WEyKPgybpa3ecCjEALbyLcWJbY1
55tVvMWDjtFJDyZFeXRtAAVKbExhdcSwe7KGEWN6u8SGHTdxlZHdpdlI7f+Vy45iABrtD1bbcK08
h8q63cjlMZ56LnJ2nlK2SZXYvj+TP6Wf3LfjKvzRqq/TynIJXrsX4H14YoSc0CZjdwlkNqHImx5c
83rIOTg3rX6VrWKTCwBmbu6waFTWNWfr1RfeUk6FyEPTpw9pGsNoHotD5aq/gWy2OdIo3j/g54/d
mJYU4ksjVidSqONn20VQLu98EfXZmMTbl7fiXw96VOb7f6P0YMOUeEJdNG9dl+V7nQDNozco2BqU
SPIP0jNPve0UDhrINoJ+KChvy0f37WKOy+9q49T1dsvwMEsFMeP4HudjOaX6YaTWAqZAkt0m6NjP
HRD8UFdZ61Qh7LUW+D2caMK1iJJTsgleoaqNSGYmKWskss4i7e00ZsIahkbywp5ty1gGIsl06zIi
tHM0CxHqmkO8gUUhJlfKpKe0CLJd2Ypk5nST8BE8azE8ap7pqOE2myqLU4FNRmOpO/y1ZEu3TdPE
fEeEMt6St9RZhRhWWM5uvOQsIHqSm/kFTUXcV1HcRRFnoYtrdfof2fzSjzAsY0IyDC96p5SJZ6Am
dml54F4vzxE67yeFd8kTJO19L81fNSiCYF25KOeoHjtTiHBs6+LeBpZHusAdTFYb0ngYvTa0R349
NXNfGuzIRLA+GMFGhtOE2OTD4K6ndHeYO4W4BppWXK6bXPb9qJ+fl5+gldb6YTN5L8NC2+75uj9o
D6+opQY2FEDV4V0pKWjHqK+yfKElSD+kRdELPgCF6pWqVpOFm83kAM4oVWnY90afIVrkxqekDz0o
jEjiXa27bHTVdyYNjsTBbwc5MQgyuY6SoLq5hS/fuoF0l1LtBtpxMWNBga+RfvWeNw9F88BEcMX4
3C82bIhpY0redAu4ObNiDvbMG3Eo2qqftoa2fPnYTV2XfHJWfjDnT5Ba8u37fnEHQWdwpgCORTPp
HtaWT2Rsw0wcVS0+KJi/Qiltla5nal74Hy8o+cyg1B7ddIvi3TOUyfVvi2gmGjIf75z+B6MW7cy2
Qlx331+kTbCcEsixswSwaXzOsPZuvREhieoquin52UCF63FY5965FztWfa0mWl43n+CHxsBREkBs
MaMcmg3GpOYVOHxCD1kmDFLhF48kVf+s0e3wlxjf8mLw3qFosH7PN+HjS6XbTcnGFFNfGeIZja+3
ulKZkdE17mqmL+kc9rMfnw147pUt0N5bOgllfy/OfPxOJqh+f1SQmOuTO1L+SZdXK6jsr/Ecdd3r
VxlPL5kDgIGmBwQrcf8LiYU5FCMVN/HBtPKBWDz4sQ08quKG7dq70//FTnFSIpaoLRqEuOlplVFI
3TAyOPWY4PmRs139ajagDZ8E68lMvthHb/VTQ8l/TZ0jfyCAcsOj9R+2DwWFUUWsn4jkmhpyyibm
7uoVzmoA0wSQIw6BRdc7F65iuy+8PfYMLC8zvnuD8QtfybDcJhr5Rc2rENOKtsuC6h0t09WNGy74
pkajOvG3Dw9HXAAO0xdtjIJcn/LDCLJgUsTuO5JNu4Fv/0h2bRcfKh6SpLzF8b88Em1rZpwzDb0d
7zW561Iqe+f7j+jgeA7kkLY7pe5RRGM5HflqTEotIuW+5beukCxl0a4WqKu52OCd5qeWCzCoPNFU
am6f5m9dxSzqm0hxL9b8/PBBlAPi8CaRpzxDv9WNJzJNIWjA0CgQWwfoGPTVL/LkejXtWgclUfaC
V4LhFhALagKjsiXSo1z3HBjyFFU0AY6X5o5BoChn1eJsuhsPnkk8qA/efxDpwq/zXaPw/hCFXLsz
rby6DHDCkZ33sS2lkrZeSPwp7QH9vsv/OGrC1eNOVy5FZn3VEq8lGMIqL76S9SOyBfz0ccAU07Qz
fDtdiR543sgIhAOU21Ef52q+a8+Iv9IeBqCYbpGIAmdIUUQT9zhfZ/VuJ2mmbQTFwz662rEtxfOj
Feuj9+q7JqpG2iqdI0pMVS1iaSOHSe6f0LQK/EG7qelehkPGlq5P3YOU4qNNAE3qAYzwH3PChcz+
d6re1HF4M+WEHPIMz50W+VvhNQrv7oPhT5lvgD8bxF9ugZSXAP2Rl1/FKr14pZqWZ1obY/veWMLh
LvEAoB4ui6XWEyP04Qw8L8zfCJL4/5+D5t2qEW0NySB3lMn1bwOIkR4qz1YFSsTIcG49LI3Nz7NX
tGWhQgvzrtxukgEZTezpGKwh28rBc96etdS8vmfqM652DdL94OnzWQPa4jvDhZNZ0fxdggMxQxV3
LeDflEg8Wm2gcfkxfCcgpKRcsK5ODJBb5JInglAgmdhQ2rsDQW2EkU+ouZOsyVEqV7KnSzpdGKe3
6gz5yHaRt8mAEotnUP23r44iPMJXZ2y0n6rVQblG9PpRyGDh0MwlMEI7aNjkuZKXlGE7NAsEib6a
pxHHdulz8Spm1GCiDFxorIs5hg6KRH6hC5o6u/P3a+NiMRqPIHssC9RLiJeTwq9ZWhcSsRI5B1cT
fnhLErngYWp2RniB6PpDpBEw2Z0fOCz9LZHFNKnLyXoaQOp8HDLzFpV6IF1d6cOY+JR99P/It3HX
w3sua6ceOng+JWUUtBRzrO1FO1GpMeJHeszUTjz8hZBvM22FHJdRSp3wucNj36AheciLgaqYbmvS
wXGPV0+HrWG0S1RKow5LltvFkPNt7QD2qZAwliw8o/rUHi7fLSvw8+vYGn38RLeEq8q+0fo/kUHx
v7MJStPEN9U69+kV3veu4o0zhqTf7ZiMbwlzt17gi1LrwlArJxNc0tzUFOLXBgeA787PYGn1Zu5I
mtMRSailljk5w3ZUeSHdiIieLM9pSI4DprUtWfwPA1Ckdt0alvtZdTyyON3PyKAlQx5LmkfFfclH
c3hWqtz8zqag+ceQKdBtwO4p1o8T5RvxCtR0R1iuOdv4cxaxhAVDOH3ioBlhDA9v797Rv7vEV2O6
/3c8j9xbHa2gUHwwyR4W9KhrzWG6H9wrVBD/9AnxANcimu4an4NgsUmdxPxpgIJwhYYEEDWpx3Uc
1ses7bStKJIbthTbwFQBfg44vM2nO2jWKOsRy2swkW0J1iotG0kx/222z3TWYNw3OuTjjY5c1khu
76pfgvaIFDOSSAcsKeSfpJIRfImiDozPEK91uFSrXpehTpPat6pAM7G238LeClC54Zdn11H1bf48
I32lG9GkRYwAx30fAUXAucT5U4J2vQpWpo4dGhZlLbVmjnAkCzVRHE+16Q1/gkXcrZuSRxYWdHf2
Hpy24j2h+dvJdvnXZHJWeQOIBR0vKYkkKRWcxvOzDSeujLYknB4OlWQe0+3HfaAKQkX82GPiAtKy
WgNFhw2NqpDrjz4tewz0qQt4e3iuN0/BJR2CyMOxjHscd49zr5tT3L3Zz5N000kOCtDfoW2zqq13
lms1HLqmMBpoPp4Y2ucBvauCjq805Zv1yjPlznQIic9zQ6KdtuAmC7iwy1Z9sTPog50aPG+Rnjad
wAZ6YZLk28hCP0tS+veymhSx2687tW2QZnGzFeaBFti3Y3PsyO2I2wqQTCznfmtlSyBlE+chk6nV
hHZnNb6y7eXyKvKG3HlRe12nabPw35fhLL3Nij+/bJQ+yWoXfwJ1kGEJ2AwF2UqcQDOvYH1n7yDx
9v9UVMwEpEk9VA5tlIaIffrW6ZG2Zf4haZIkhKA2GFv7RN3yCl723vL7iOZPeE/SAjfRLv9ckJww
iDJ8JsMZdPo//vivBMRWBXkLAvM39v4xhACO1pyt0aEAp14na+e0Rgx5Y7nrhQSWa0hhNCH1i06d
RbfbnK9QcpuX0wYUCcH+tnYbGcbl6sN7aeYC5kH4YX5fCAUJyCepBbpGddHBbAf4Dj2HxSDeB49e
JPoS77gwfqr8M5wGMZpkyuOcR8t3xWUFcRbL/LGSiVsffHN+Dsw06jRH/SFofy3gLpNOmWdbKXpi
f00AdJ9OEr8U8Nx4l9L31kAXDuKAr0ZPaRZ8q2JfZWEc9dPMzmgRET3QfHIqJrIvLf4AyktGxwqC
wuFgEZQ6Yk43PDudvg5TECWq1ZOJeh+QaWW2btPmk5KM8vmyoPaRbTHTyKbcywsbahUsx1a2dAUv
1wyjZW4M6CmvmaywGur9JEIlIv6bToFZLWuWJuxAAQCnBuYnyi9NiVWM8JGmU9s3w9JiH5dTHZNb
tf2QDy3WIGmj/pMqzXfc0ZGgzyV7EVTyiKRSJvPXjI2V6VNm5/4P4t5g7zMZfc3woNN8ZAhvq+zi
StuEqgCCDRaLTaPPkLSc56d5fN6XHB7zjiskyx7wnEfU/qj4AsRYtqjQFgZgCw2nAMfYYZ7oEC96
F+5PISD2J7CqdQWL/ehhS+RgKAvHKrQ7hy8wAuW9E23UcP0pXNwVPTuD0p1x2DKnLv0axnGYAWFW
2qymv0ilKejyzYBadZjlY1rLTtX2shxXBGt0mQzhv9aTTB+LlsAc3FMPzW16cN5/Tdt/VKadIAlQ
2PYQFVtCkgEiQlIJ4Aygt6M4Z1RgHlMyfZtI2yWwBkHJ7QYZBVQD2194LxlFcU5Z0CnxbSdLZB3f
YEZYTUBvNWl7DEnbQclSop4FV/0O/vddkFxtrFogvoCVY8NRoapE72Njmd1Fo1zUjQWvNeMb23CT
Np3QiSFeoCFdVemtVq8cCm9sJ/hdnp3Z/7ZpQPb4DGk5OJ2wtipXQth3idx6b4bPt1tUU7KPipzU
lLFoxwiPcaRh1g6qYCGtU86A0vJWKp31rxBAUK+//OseHaSbFTHyOfHU6UDRLEy5VdXKnbAsD2Fo
35KF+o90sEW5zjsnR3TwS6OLaIOgVJvIEBZZgUDNuRblHDx0+zW9WlLNTiIbvAx5COrqdpqvsHCf
zpFV+aGuTAPLcDMUrAxpWdiLlKOPu1Cgxnx6+NgYlPbGSmx6uBusflQpFStHSm3z/acfG4j8bIYy
5PYR/jost4PqNugCwD/lkmK2VrI3TpS7Oju3a0zw1lEo1Rwk4iK0prFQ+LyIkAZutZACYaxYGc0x
wktOAElgSlHZNsRh9NtnXynEPxEbqAY1I3B4ZBXKyBjrxgfAns67OI4O/yjYMeauJl8HAhgn6eft
HsASnYB1EwLItczOozxpVYQ3GwCLRbgeihUC/VKbezDbjAblauf5prEWOpeOekNWUU1Sn2v1pZlw
IG6avZSxtv30c6bOabpVX9bgENyhhjnqlD3oB3Q2K4Pa5rzmw1t8uKI6tmMSMayUPES+VG+37CWB
NhcnmCS402sgcZntzMjLLekJszhRn7WhW5OYO2pcy9yGoNk8cTKeUtNt+rB+QvaqCqxphPc66R+1
TerSyhSe731PB+sAOGHDY0GORnDAoZbl25OkOF4JBk9LN/ipxR4nhXQDByBrh05Gikq29yNyit5w
y+ytw5ajgcl08sh6YoZolONu0O6yK0v/UTeGGsZ/6r3AVUTNq7wt8nTuMJzdY1v8GZ+bLTzgfCAu
wUlgfwagkQNQAMgiUz9jCXYB2uh/SFh//clGFRyCCK4Jrs2hHNC3WjLt8t0X0Ie9R9jqmGX6WylG
Rue7A+npUKRohNozT1DievsMAZ52enpp1Vx/BOvF1YbJUmmD0dQdfDj/Us814OeDQEjlOhzGcKCg
KBv8kRosgz/sYAjHbUV24XiFs31piRheod1RP9CT6O/fmK8YlGJv0a8QcgRDrE6LbL8djxlhiwar
NbCsZd5k5YYe7+nB/0BSuvJJWh5CB2Q/xTiSDS1AHwRGa1pJyLPP/OHzeKK7hcU2IQnFqzGRQuZM
w9L316tnErhEbONQj+KJn9jg6jMPmO471i77B/GRHQFpPzCKP7vMgYg1Ko64BFtKXlExMmeJGHo6
esEa+gB0b2kLoRRhfMInP3A57cxlZy2qk3Hdgy2UsK/Sv9zxRCGW+bm0ugZhY9aL8gdw0ILl/nev
qDV31Mwpj6xFloPHwWKLjZ8Tw+Q8JXTGRMj7HqkKbgGAv0sST+fzcvDIEsEtO8qAYiWB3eEH03kT
pbh2951xmBvw1gIOT46SbOKtqd/f0u3MBfUnpS+e+0JzuE8kFzoWImIYdVkrvGAst03W+qAMxbMM
WLfUwh9rUG5UxsUQjNO3Fj0Gu+5B0elCcK2B+fL7KRJ7tfNy44xfmrMQkU/rRqamgn9TeVmBj0vS
QRfXcbg82N2nW8VXoQYh4vUreep2D3iP7MKlgtfCiME6hGsRMcx9FtNhe7LilZf7dgS7OExQ0lgc
Kdki3vVbKC1pqwO2UXzq7WTTB4GY81Cqvvc1v5aRbuXiZ7ApCIpRrx99pKNGXBT/3cfHNX8Ks7Bv
nAadO+Uu1RMvJXIyI3UQxrnYruqVrrciQOtFjigA1GvI6JHz0Dnqkqqcf6pEIybipo46jgayyAxi
vfIWcKE6LA5+P0kXKz0fDEjxRnPJytnt2F2j1tJSwC+0ZlCSN5+ONrgjZx6Ohj3nz5jKmfQDgFUb
jf9fFIMoUmSpxQ+4askSnJOfrl0ffC3RnluiCh93MxMZxwosRa8xL3J9p4W3wtdBXEA8yqWGvF9I
KgNpEFLs9M+6Rs3NkizkofD7+pQKbc6ZEoh3vrWGsyeNDxfhDlAaPfDDymdRkBSc2FI06snLzaBm
Lh+1klD/yWkVDt5rTOiqfaKQNMWVQjJ5x+wFRwnIPANxUg2RjGKdplowZyek7z/Qw8lyxb9Ebhen
ciRZLMIJvpmeKO6rz517fA6iUXzM0bwJrpeeoWi6RI3WxeycmwQLX0UpNtd6gGqblBAd7jqn/DID
SASbm21+f3VSC+MV3FwLrGjua2/czYOKes6iJcR64elvD2CXyRmzt+qn3d9iHMBlNZdzV3sNMwLl
0CFFAHgu+wDclpxboBl1ybQRPKvJjdOf1AqzUOPRJ6IM+hkzWOLJCzp3W6FXbwFXtJdfkywXKWAW
q/1bttFPg10vVshW1udy58gpwANQpNOl1X+eFJJ6xklEtcznfadTFUYkccMatVOdES5c/nONhuJ2
kEW4RgP7DhxL2nPUst9+4Ai0/ga+kbqqr9N9JU+/U731eU/g/uCBe/uIxuR2tit9QfjmHW7IyMGM
qJ7DccmQCrl9ojgiwN9BbOl1PtqL2IWIu2NDqPd7+Xj9B0oiIl9M3F7oDQ8H6AAO38D32AMUna+V
D1yrq+4JLwgJ2b5AICJruSCQH8SvrNrgt6LPFS99q5GIDYwY4VK1YP/EDiDAKJJkLr5gQRgl4Kpv
R/0xXqYDaWrGB6Y/byBIftEfKXaI3SGcJq4kIbgcXnVYFSCFpmmlaW1pqc6Df+jqTBso4mXmYzPp
KLAsQAUr3qPnLeeif37XI2Y6Z9HNFnPeKU0EA+6OClOBZ+CPHWpFv38k2rVHPotzWnmnD5iy5A/2
IriiwWzaQQtmInE34GSqBmwX8cOaOktFzHrh5xkrmdMQjRF+hb4LwTkXykNb0fg09g/S6sVVN4CV
ANgpvP1ZrgFe3/MGUK9h1Hdheab2FiWdUSV8B8/Of0rj/rLtvJbM2xYE81kIcba0f6FiIDUQ55fd
pb6WpTgwn9/WlV25/dm1yqVx3eZY3eOpb4bcbda2Dr6ziMflBPVKKR20VAatvtfWAltQYblf70lF
5raz46wIpuepktc0G/bTH9WFe0WG3srVWCN4nug2j7qwh4dPjQTCoSrGSt2ksqJQwxrG+Wm23i/x
RlZ1xgaGjOH75AxfmaQiEPpAcqxVG08zNJUVFnRbsXTiI6PDxT1HP9K9rr9h26f5dgO7tMmZ9Kfq
KO8lzOGrkjUndsCqNSWFms/9tKfKYJJdC396LizObIwcqvV4UbQxKpKC45ebvcR59wwsioX3qUYv
uKbtzspCeQx8CPyf8cjnzlVzOpFtTnx4BMcMtJVnZ+5++7u3q8bPzoGDJOpEvv+mLfWKU7X4OnU8
P32f6+L9Q507dMduuOCUAd5dT8RNgGa2AhSdTCpFGd24NER3IC0kAnUuc2EHfJ1S7Apdv0LHuHPA
ClchT16IE1vuGje0wyo/DZO9wVOIVn8q6uxLsjG0sRIgPFRA0G0vFsAiGfepTP1cFuYnTS3Uyc8i
WsK1+XQmOtiAIPuzIVS2xIROd6I+H03pABfRbhgtIgt14/fDd/IJUi19fAYe3JrQFQ3g0IWJdCVK
ecDFpi2YURxpttEbeZtTJx92i9EXTUoYakMDSpMRzT2qMdRh5y4dy2uYN4mHby/L1gkXhcbYv7yD
TptsvwQoXMg7Cviaggj3AlgfQcYC6fhSoUgR5GupQDN+8lyZ3R1nEfGTrP1YPl/vST+nkHkR5HkE
JH8jTst+n34IdGP7kR1P0sA2t6gZeR27AXqWhKVVgV5RXxuXQVO4p+a29s0FJIAG2aM2Pi1ugMCw
2g55HbZF7rwZgOGtfDpf+yAW+egQHoNgqVxoDwREto9xKmRkklPXnARQpwT4NKcIwRVMTa04lHzN
vw7n5VoKm/kBuTtsafxpKZquLsIR7b/BzpC8USRujxIBQKTh60W6Dr9jT7f2lcW9K/Y7n56p/ul4
3uWxbXwziwOQn9DtXZp1sep7couDOe1MMDL9De5qoeYQpVCa068e+ugWTogjyzbhoTjYs+ToFS7S
xwtDmauv4uhx+x7ipEHfjCn1162ASiSm18e/RXdCW3dG03jZZwbbrHxnAC45cEvpWS8D/VvRRQRk
zfFbR82BPT5JMbLDxpB1dMCdPnsNsDTzrwDOXooLtL5+12zzBqMmzbKBVPKl85YAP1bWhO4m212q
Atks6LzA9RzhB/+FElzTHFiv4AgtSe6eWvAQ3rw7MtHnQMYUfVHcAaiGBm99zCMQsfQMm6TulG4+
swicOwo8pM+a4t5WP9aA5qFV7A5+r2D6cgPsH9UefxVLlIYYDY6Bm40voH9RtK8WfxojgIGTRMTN
UHzSF/xp22wmWqzlnM5znpgkToITV85go7u5oxPJga9NTMJt8mQxg3VmtEaKFpQ+PmdJ9JzrRCY5
r5HaUyQw/LX5dthXAPI68Wz4RjrOKqzkP/kfb1CQ0uEdhpdMtKjsw+ydg0iTYVeisqB40do9TMuu
cmuxkZ95VaPWQSFoe9Xc1FxQzmnXc8PXG9bAlOaba6ZUbfziSqJppg0caE8elF/ZxrAdTMQjgwMX
F/xBhqcoC6j0vUrwor1hAamNAV6bENl0a69HKAdLkA74Wq3R3hs3wNHZ7qtYn9HB7RUMlSn9iPd2
hUZHhvXPZI7wrTojeeILubICGziqfUwOIHc44NwwpEGBHp7POYqDfRQgJYdngxDZon7S24rio3PI
0CMSBPdV6DbeKhrSDBgpBvWhrpzarjbipD8tbg8JQ20yPrYGlV7XQjEUWAmmAn4haxrnEsDKFV8F
o+XQY2z15IHnyQkVnjgdpM7XDt0Sq8GNErm0hSpUoZz6mqfIFbdFcWh4TSgpYgwQajEmzNr1yj41
x/YW8vDgAmzs8Gu55Wvu4Av+JL1a17Y2E4wt53iZQjv9iqIqsMASg4uwoPdXEkm+qyqTx/nMCEjO
Vy3CjgpE9gItFKdpu3+t2ni3+eAd4GWuZOSnR717erCWvpvuMdci3I4o1sHjsnPlV1fj9F6Jlqwj
a+j0gHfSnmrsijSwbEr8PlwshnlG+KHSm4et8qjmyFomiAA63eK5xzTszgzRQ5Fph6Sel6QgSD3Z
LUu+FZ3QwmPefYVpH5fa+6lV5w/HRkO1JlkjKBQDHus2UrDFIZvyOUPWIK1BM8tab67jmahtt2OG
99U6m8btWy5KF8cFZoFS729v7rszAF5wcvVLFGUOL+HtDztb0aMOWQn9mRm6cZl8Q5oRxPUPSrdp
wC2HKgAE8rgxXBFnaO9DZ0nM/GvTGS2YLrKX+4ht2Nqnnqw7IeVxnoZp+Z4xMR83tN9xS3OOXhnt
0rhyDdWXdbajWE3XFZoxbmacadMM6OsRizRg4m93oVvSQsXFdXciK632fVd+nmN24jmpsokQ5hWs
ZzE+wbCKexbP5WaGAYEfHs7Tzq70uXOUWMgGUJYnMhiS9l2OlF9oW6ryk2+hIe/ZDet7vDQlQlVI
+z5SW/Xx6pLW6B//Av3KgEvrWqOtkzUyVFsV17VhqvP2xsPO5eE76sKta0dV1ThsHAwBzTyG8uyn
dHToD6p31ZB0g1CPajw9VQxMdMTR2WN9Yx8xmIglKY5mbZ4ws8Z7qzoaB1EZ7BOXufDsARADXUIB
JgcZQS3yvyYUmQkPS8oMejz2B2mf4Zy996coXcGieo30Q9S/bG4tqoGoInzBmVvgzt7hT0xvIVMu
k9Rx3uU9DA7muEC+1Dr2hkLJB2757QWu7Pq9KjovR1WbhaAWDDLFgBGuWZ4Jrw6+CizkoKNlEVRF
Ur1pq1tiEHz4XQg2zoeoTrCki+jBLN3qs+tO9ha2Hmr9tx2eFCaSGhWOtzTfBZlhF1HcrawTZUvO
231bJvTGWc34tiLpJdz/phQYuYv+iB8OrZz3AanuMvaqUKDVOHV6OI4xJ4/+cyXR3IQ+X5Ukov5L
/bos9TAFCW1GycoiWAiL+5Rtn6qRBBgvmCB0Iqd7GMP66cJf5S2/8fn3eU8pDdziOIMKXDNjqKi/
exZu4WHurdKakxqUefJBlJHOGM0FTSFVXvKEBADQxu75+cYp0lrGRaTj/mlHK2S34JcQkS7AYVVy
PQOVlh/S3eJJ2cfqkDvhFcK/SccU2LbUJmevdSVF7bXDlvFY2G/lw06jqb9ChWj7IvZu5S2kg+Rd
+1B79JfAHRoKICufJMpzXZmmNcNMZHgBJwLyFOHeAwynuV28PeCUC3G122jrNo5NQPKa2IFbo9T9
hlHYgFdPrCo4lZVg2f9/qfkVlOs1OFML78icazBOegNRjpH1jsYHe4/PiIOqveEXP7nqxGyLuHY3
Jdsvj1LG0XgMnJmJgVEHaiPzjkrGQ8kfxF0I7ahSb+MCBiDHBNLm4KU2Z1gQvETe2AXa3BKIVM7i
gRgAJi05lMTRn0yLcHmIAf5p2W1oeOqAcCQ9myHV2T9cwzNklMW4yB+htFtrUHvR2EFezSyx1Wzu
YnG7dQ0pWOYuejOJ9KuwfMY1HoT2xQU2ROvN10nRo1jGsEBWvnlq+GmFOoVlTJ6xGuyJIQSV3RJE
WkGrN69xeIdwNTR15Z6ki8dK/RrDV5FTRutYG9fXuDx82DQqc72e+0xB1KQDaXnPTW0wwSpevCNj
Rc950Yp06ynyjl67LwYUdbK2MA+JhK+8dSYqLFNaZjlV5arrzWQNDaeeknc+mfsiv2Ed6DZ/+m61
4ZEqXQnV/muCKehJ3OiNxZLqxEkVptiQo20tijXmBJ6Gb6MryahHWCwZroCDoGSVcN5bZIscm1UY
HpWD6S7PLGWxBziOkPc8r77NIXhhm5L8UreDjNLE6sQpsyf5PBGBYm7aMXp7L5LvXVYgnAEJBJU4
r6fyMelELmCkLd/9vFepotIhpjtAqOR8u8Kp/gcxhDWZFxXzD12opaZpFEs21jAKLuANfjQaSruj
nJS7HixClvM4ken94QJEc0KDqedvHaWYNLfgOJH98u6tMdYUXEaO+4dYwFD1VnhBBMIhwX+znKyq
DMGh+8SaouTu5rTSORNW2sFi9msDNgo3DPqPcspVosl1OffjrlzU2RQdjaN+rM2IFSTV8BsJxWtI
+zAU3wSchKrXIUmu+VxLKaOv7rXq86Tj3eZ9jzt/fHS79EV1Q1SalDabRfh+YRFPaAydhNOczJ95
Uk93rl7bzglaJf+jRYWJILcqr7NzxkrPEGTdK5sN8c/aVJ98Gc7Urd4CmgxOHahXqEJxaXB8CtKJ
ZC/IggLjKrr9uJJDct6htKfXqzkfWDfb7QZwB7j8zYF7KZiifJkOfwbfrkOTMCeh8Tv2hSQs6W6Q
Fgpn3Lxtb0cjyqJSs9d0h7cRAhPya4GRtbHr7/TQ7b2M+0y0OlmSYh/GOdyXN5zKTT547njlw5jw
PkSMfHafuT0E6hfk0No1ho691mjbnByo89Zem+BFJtf/zZGadlGOW5P/f7WSTnn6YdwQpSBxbGlZ
FVuHxaOL4ip6DaaNUbREKIDXR9k6ezM6+DrRnvCyYf6ZMTtOsA/KRBi6DMGerhGf1SQP321cCbTW
3R2s3Xkird0qFBpJDFnWIt1UO9XUaMI1Ti/AiqA18484oBeKSjXG9mx0r/uLTA+bJ+kQcMmW1ivr
qzKt9aTs5raD/fmHztixTfbuMLSiiyDbNSNZDNqYWqEJjDwH23Y6utRlwOh9GqrtcIOaw0veyMh+
8vh9bGTWGizliR2B7OI4STd2M9OacRW/dyMLSLXKRSTNSFGBM6J51399YnVYDop56CZQBDGKgWjd
w5uWuZ3UC6aGPL0RJoUBG+SccB4Ndpxl2T0yZwDoMgMd2nPyOUx8jZsV1Iw/cOtkGc0GqPC5wylQ
FZBqLg4OVeACLh/ukEVOJVXcrTW4x4LbugN59bU7kXs5LkNcYs1wLqyqOlzEPYyE/oyaDdB9Aw5i
vND7wOSidA25IPgpUx1GJKL9fZjqxuKaSLguwF1i32ib00502m7dtS1Yi1cldugvcrZwvFKxX3BQ
Vy+9mVUh9bfb5Tb6t0kk4vafZqCOuHOy1vcLpqqmQY8E7CDrzm3bPBSpr16oii35dCOoeeyQZQiK
50J05J6sLQvA3zp8gy75QXak6Sv93bJ0aVEPBCsgJIQEWnc/jSWTy+mDoiEnCxcNvz6Dik8op7E6
sVVXprF1wweI0bmbQcW0XBeEHhiCnZEzS0GZPjbH7FFRetV5LeDhl3RsP9s2/op8mDFwpIFybx6l
MpE39PFSqikr1NT7aaBG5rQQHcJFqzXnhCQlq3+KeJRyg2QwgIul2uG79CcMF4eip9VwUe5PNXWq
n1bA3RAq6RXGwkT1w8WiuiwWaRaHOmeMCAekkkRwwfkEhG078HUk3UUaDGCaAz89Y1m+1VwBlNY3
XzKfMGJ/HBbJjHrFVTshdDw8MlgRAbD0aFXopC//cB3qDGmT6zYpTscXTZ8G7MBkSgSKXcTnMceh
tIITBDs1iZQyfol96d2Iu6ezS56mdqWce67RCK5u9UjUVaa52spWI56ZBB9mRE6Q/Nw4AJhSKWTM
dmLR4lf71FtkU8aHKdEf3M/S6djLKoHY8E2DgMXLJqLVq2MU5pLySVQc1xjlIbZhjUPWN21B5kj5
9RyVZneywxBdeBo9fAn6hf4v5Mo8vcqDI9NQpI0W544mJ0RdK+QliN306SVywpBXFUuikvD9NUJN
go9iCV/jngv3kZcQ8dPsKeHuox4mlM1fNiSwpUfL5KqkeoTN2N7DCQD0B20s5XLIEj7B8UnnCDOt
6MaphxxZvkDF9aKkpdxjjpupHj2mJtEbwDDn253KAG5aF47GL/yjklzxylCrDPICTYTNQjSu14f5
BCkuFEKFl4a+k+w6AyzVmMsaDjXkwsJ3a4NhdsbdFR4WUgVs7p9+KIVoYmChjbmoH5YaDQoG93xl
TfCYp69OWhqs9rCpll6roZ/jxJJsoTHSAEHcFRam3SZkfaOzmY9oRQaatj3cO/2J9DUK+lxTbPn9
6E54bDbRukQf6xuuQRHrM1G3PjFASdW5SJDZUIvDRPNVkW8LyzRG5NQ6KHnOBVQWjf/vlAfhFEnq
l9SjfDNaoycSxh3TftTVDhDvRhZB1ZsvjoNU2wijy7+BO93+FcMiXNRHb+N0EVeb/juCjG4AvUU9
E78CH2ZtO0IQ94YHoM7SgdeoTTAn9iuHQ51BO7zPn9qiK/dK6SqAQNyJfu0syMXI+wyikH/jTfgV
ntd7Ri8U7P7jekhEDkJieZz1Eb5k1MZyjUS2OM9+oH6cJd0xqb8r7zlnUw8ZR6IFcsnbELYHkBId
r36IFMO2bZmvTKNYqebTQ9cPph60YpomDKmIvYBgYnXg0Z5tQY2w2ykGxalI3TU/1b9fukSQP6u8
6bfR3ic0maRMvWTp+SzsHt4h3XJg2pGRsh28RkmxpfVRVpoFq3exAlaRzTMIZrrsQYaXzDsoNS+h
1C736+o6Ua2GIBMnWjOIXaXl0E6EXRr7eCM2DFe2QT2eK1/AKJ2kFLhqczBAhjGxXb3yPEh5+g/C
2kps/071yjJ1hYBFf5BUzSdyFKcQipaULKJMx4valP/Cy30uOS618y+BzIzis2JYpt5xkksii9Qx
VWQtLWAsg4jz/+T+AFKy6sn+RKaUOBu2CIoVNrY1VAEJsgaAKP4+P9VEZV49CC5VVhDrkoTLs6aG
aH66GzxKL95KDgFOfgxc9TpFCm6ubLkTnIrO5Sm4G9fqnb9MEKi/kyhEh/25osvEvK3PgtYt55VB
bKBpCdWLivQIUiTGa0aZxoVrNUivet8typimhejTV7MVHlt+hVhwpaDdA5N36GGRbH7V6y9sZKAH
GVaflaDbc4Wl3+7WWdaDYlVnSCwLSlNPAUcgiPw0q7Vs7U3BphTTVCP/t9KOf6MRo6XoGz12ILjk
129ZuO+Gsfsvrhi6nUCFg8fVlkQ+HbTuld2UCwmd/6SX3LY+o0TJRojmahZMizFwEZInpXyGOm7P
DWCGQm5LsbsfjqqAsFX1q9lnoLBtR0Ts1tQRCnFbgR35HesWrNWqUWr18rg86iHY81zfWSbTcXVB
ZYjOsK0rohD7DCRSDAoZeGQgtfWB+cIUg0BulFhCTxcoNjfBFw8dtCAYYsf5xp+jnR2QzUjYdNE2
te4UHUsYHGU9wIkhCQQJiUj2y8jCbnT5NsNWkpONl8KbNC77YZuRW9PlS8cD4dFQNRBDEkSqnb1w
DVljbOiVTGv33Lww+LqGx2byWGl/fTZV9yq2FnjeW8gjidfQbRbgQb8vdswNzTNfZJKOhXHFWBQS
vSfeTViOOEFvwsChT69R+ql0iqlCnL34GGPX04N8ishPYZNw6snqxmmoCuLQFjjLmz1dEy68xMhA
MRokUPDk6enP7RWqfPjJgmXnImVwicjoutOd6GdECaS3Nh7F97kGgtnsXfam8fLPI2gTz+YRkAx6
SS7VnoSl5jzM7PD8gYSf++nbNFhyx/5ChAmo/1lM2JQGcqo7t18FiXyMmsFXgjJmA5EQ2x5fFjcD
4EOMU9LSZotIYo+yG7l6rSg/8URzuxTkKxu9S4/p6caLPFoaYiE+Dhy9RaoovBa0imVR1bVjmlJw
AWvu8MHf7BcShonXispvkX/yqdNaDqcIJR3vgmrK/xOU+n8ZXDaFX6apUr2nVJhVMWQdtOKeyINV
s5JJoH6/K5Wvo0bZUQJiBSJCjCpTPe/gUHWrxlaj/AqhfwY1EU2T7P2DMXYxoyNX8306m3FcCihp
fIdNuZgfufJamWaVCVcN/pKpt82/aovC5CDME1hKSEyh9+7SGKTFnxj1D/8w7/5Zk0e0fO6+VWfU
USSFgC0tj7I5/+iNIpv6DFnZUDXjHef15PosBx5BmWa9WY6NLok8ZTNvPsBjKDIPCzuEwxINDw4y
LYuuZIB9n3OWsu09hd/OVB1lhELQ7YQaxN99v/80FBJePMJFscB6qc+XlxvpEJ8zkAvB259rdBIu
8f0cPxtKHH6Klo1GCbV3Ai1RREjV+DK8KNMVgUNuSE8/amzUsexeCPU3lfCu3Elmvj4luvX4WFxq
v/4Ra0XgJsensIFgc+tSM6cZ/gtcnl3i5rJvXt4hbpMy/eCej1cKOuI4C3Zd+WMCsleNiHIPcGBr
9RS3y6atwlykqO6kzPnLMbn+viIILyqfG7mlo/LNyl7JzmtlHwoR0RZ5+CUMF51Ps4yMVGzGr2/E
q80q7r1NBnYXVEWv+E7/mwYhp0dgQ3I3vjvSqQ1vZJPh46GiCq9Exde6e13VMT/5KF5s5NU0yN8E
tJFMAHj1piGb957tNy5OvUSEarOr+CydnNovoPirR9I5M2ockqqY6P8uqgYT9dstlwiWo9O/s5zU
LSrUdMEyNu6Cg7AT+FTpqBv50xKhqW+qS+32EQ4/Tm7lxo6ZIOjq2Cw6WdMIhcY7aRS9pllq3iLg
bxjA9g2gxQ9+/Hs6TXVxI9C/eM3dcAB7FvwUmGUhZEmAZeaHr4Q2W6736WKRi1PTX7sQz8gKMX+f
bmuA5kiceHcfPTNM8E7UUOfPNyP3o9k0h8gspeiKUFM9tOyqcavLW0tg54KTy5ZXNo/fRkX6+bzl
92ZIAZqnRPrUxDX+Ae9Nx/w4fhqw1SRFzReOIAHTWxgsIDJEQJon4/Ytt9gtpApTkyS2/MjlTVL4
FnfwY7m8WMA+OcAVBU3T0m+Byhq+xmOwVay9RuVTqx0QA4cVZLRSyFrngqy+M/bWkOopI0nh+UtJ
4RdiCMymNAxZ8DQP3a1Z+gCZEmPsaeSBBqvaBrsRxy1bdVk6iLJk1H1ioxZUciMVW2jHIWOu9WcW
uuoUwWON3t/Fs04lWwiCigsVGf8Tlc7dAE/EZuA8fIH7e11nGPVnoNd/EBGKdKH5ATS14f4vbGJC
P5sdSomYbXf0VqzxXBpVbNBbg9utqBl3cvHyezrnaMYYZcjKBkqVAZ2jpFH8hXLNHieIt2HoGuYA
eTbP0d2jxziV1OuBuZ+9T2hL+Rjdh9cTYoscA5EEfRLm7f6msBkpYIqEbM93Ws/YvrvJEjxBblaQ
JwVLlIEsBKD8FHeTu7/DAAgtDXLnJovejEaOdSGLg5lcqLecw4xqEOLiiHfrTNCbqCC1rxTUSNqo
PbfOA378dLbetmNmi/FnajKcR7rLTWv1yb77v5mHUntOY/Nua+kEi7qd1bJcQZrcMd+VEW9yaLBR
L6sasg3n4fuMgl+FJPzTAt1kioCkIpfTOZfV/acQCuaKzN2GU02POL/PMGOYYA9Vhv/MSRGM6Wki
9IX6IEx9dyU20IVStgFCBrIC0FjhLcd93KZLMHqScC+l7Rtr3//O9IkZFRAVbni+9TWeXlKXkpdh
KlGUBW3xBmypSnSJ2jOug2BuhtSvv7tc+pFJJjlTQxy5SxKSgm6m8yJvHNjnxn/NhYi8bOjeWW4C
YOndVeY0gv92+uFlf6q75ajexsaS1dhbPv64RB9IUxYbb/RVDUfUEWdR1i/x8L9sRfeLUEFkT5AI
k8afcMH6/1D9JTDeRJhZK8bmjOdvKZqT3eOqD5JdQZk7mWSz5eZ6p39FIbO4UypTulugZtk+bPdD
UlZ2guGd+1TKdo23CsVXyJkvRW4PqPT+dWxSGPYJZjIO1UxT+S0OMLwoonXpsoxq/M7ZFvXLfnP4
FaiQM88NZN3pXH6wEhzrLLKiXx6yob56BSu4BPh+p0jVfI4990Ebw/braiQtirqaMzR+Di/m/fuM
ubifHpm1luuYTUYtl4Bbe1hmJVMmgWnzIwtS753yG6yZP9ZUAqAOYQJ7/oqgYY2f6f4Ps7Ij+/JW
0Z/ZWKal6X2ssZg76nsUw+wapa7tFFtbvIqXE5kwQ/C+hlgT25mY2QDwY8GMomiwJoY8tk3h5fO0
yPOG3BLoRjvgp9BVZ4Lmi0wx/KM9a1v9t3MQ6KpBwqxMpb4RoZmef69TYIATvv2N7jdaDblkrn7O
+/pRe4kHDdL/pOVfX44mHc+4OLRu4WPe3yAOaJgsyGzy5CSMVCUoDK7+LozgzHxnuszRMRTY1Zjc
Hfs9Z/UeII0GHT0D8BjDMutZw/CxHJzs7UoRVMvK7XqE8kRZxLP+9jbb7sfvUa2HjGBvvOw1Ih0r
OQLJzDwvU2/N/IQij0YNo2Vj/pZ/3ycerko33BAUQCKPfaShW35gJ1JfXqGJx3a/ozVFjmfNpkEm
VX66CMBJ/j4GIw+I+r7c6PYxMdZ6zfRGFSqP1eDcFhyz9Ti4ZjO+7awZaJJge66SLDguHv5BfnxF
9EBncw8YPQhIOqG6ptE+0YFFAKiIK49nq1GpnNv8wkEfTUkGn7RdtBe/vlrgf3GrRqUhLxqdKdiN
vIZ3UfM5a2+0krCUSVlcf1Js3sGHmwUHQ8yF24UNtJmr/7Si/jRtfTbOylLwi/tWc9nMBsBBpqah
MGOu/y4ZYF5tGDZdTMrsQ/b/aYiJGNnVsS8Y4AV1T/Aa45dsIYLjJuiSQbK4/U3+uUPWOXWP+M4B
KS40tKlLrcTP/aycDY7b7kPv0ARcsyUZoK/lrW/TMN+DSoQZuaRvPLVL0pwnvpsaonijNEt9CCGs
xgzoZyeQ4cEYMcjd+onVsB90TTsQNC57vN0sNkXllZKP+qDPtKe6wgBt1DCYexvT67/Kq6UTGkWH
hrXBXR6TAQOl3MzDKlpqs9HZwbRN0FYUNxgyyQyw9uKF7HkSe/nikXfVQqdZvBoZN8+P44X7sOys
AnsY2N1tqra5zKHPTIQ02VqFfnevFayO/jDI8DEK983fZvNjYjAyMGydD3JiVP5zY8zOnZfdythO
CPpAVyKt2bB8hxuOiYRxNhIkdYRf6sg49db2mqJR18DTUEqDUuLNJyKQ+EzqcX3woDojfLh7fqw/
7F4XN8v3YRZGHeP4KFTzuEQxb+XQQi9AUz2EBjauUmzlsdFOrO1Pnu+WeeHlX/7XoSG31NYPIkyo
iiDn9cuFwPcTI0n8i9g40jU5WjHRIhTST4yBjFkCnGCby1/22VRW5eLPV7/SyFx5MVpu5m+uFoKo
Fg8mEAavXFu+nY85xWmpWXEOrE83ro/yaUPVFGtIwZLI4ql6fyYUWPXzAmBCNmdbvqtvJMUvdgOh
S9Tyz8kSPjMBllFjKFBJeOGxkX8oCguyF/Xj9Sfg8IgiAS5prmcKA6zeerEdUsAidJt+ZcW5C+Di
R+4JUUA8JSjwSB8rJOQlkPR+JTaip22X+mdJyPFZIBCwU+8Np6xa1FT1aqVXkUqPLRMAfoeZP6Jb
gRoN5k7g1pmPnnBW3BxMxBGMAZD2Dnc3cQFbprknDZ56yNIDuyDereehB9GBYj2ZQfNm7WCyDrWd
SV+XyH7wJeLLynWM8P51Ih1ZWRPUsVgYqysbuDzS/OhaLNnSoWqv7r7bJpm11TK/wFD7Yz6HwAPe
AtbXPZWRVukAZYkwHtjiVBFhFmAgxegdHfT6JZP/fSQhw+qvovILb3Cyq0cYNMl8kyG8/HGM3BHM
H5J8CxhtKsE3xmoqVVMcpdkVGwbjpCdAV2bYVHR1puaGhuo3zWuPX8cIbqGptNVg/rjCb+VasAhB
xbhNJXga7Ps4NP2R830C/xAHkP6ioD6iwqyiHiA4Cds5WI/mU3Zo3yiylmiupu+3aer37wB4jpLd
BocboYrVcGjBaGMFRh4cgAVzrfT2i9FZ8V3ge2gq1uLD0bGCIehd3KgvqRHAoa8mRx9NpJSRJHFm
zjbcipQXsT+qJ1XYq8f9xKk5Y1qxoguq4MbvldazCXaqanbAb66u6O933gpTDgjGhSTGPvtBJdel
msZ9zHI6/Jowr3lzSth7+RwIsa73G9HL0f3rT9Znmod2gYGkZijSUS7YwQP6Ncpj5BkqDRTWWOs8
1y1ZG2D1RD8alg6pgDQ+RlQU/K8WBlgBQyEBc0Wb4S1MHknfaaB+hksd99+KAn8yQmzsjAmxaH4r
BN1Ga83vjx9rSW3qWlzb59IsoEyhRXd13FbeApKkTyTdHZVA0WCBIVXDgvC1RwyDD8TKf1u94FC0
zz1NkYDOyLxPUIp9tWK7Q48v9M6Q3MsulJ1bGT4BM5c4w4nfdqFoGNmElMAZp7siUMO39EMPxn0p
T5lvj7ZuIVD92Qd2DM+dUh/0r4Opnmj3+DTliQHQs88IdrGDeb91XU3c9JcOPdynXyKIYxMIKwSI
oO1ctZZWmvzsxaL1anG0PZhHnovOVl7wHrmbwOYtojsCC38oQ2C44Y9r7wtCshW8akHVTOm13N/0
scTa2uAkIjkcV9qfShwJOTJvN7o0Notpi5Oi5e0gmtw2BQ4T5fgkHhDYnd6E1WfHYd8wMFIZ3Zcq
4HanziZY+MNzjdpdpfW0kNJ/qkFTuYu+0hwBgefAGHMgx4mFYxlULV8h8FgPe/euOqGSYRgwB8X2
AmN2YzarsF0ouYfgFHlTPUf0B7tpO9QgggPtr4//sBiQTSjNQYY45q52I7trDA4mA/jSVopo8QOR
qXeVAn1663ncBm6IrEcnPnWM5v6XoCbPC4ryC8+1MgQG8N6v8gMowVO+8cxiBYWAMZHxNjeJ4onR
KX+kpFnn8Z5qiPXyis7UfJl7rbovEVaUwY+YdJdhCHryMQhPrn8CRcDBbe6vXvxdUurRoyMki5ww
DDOMMs9Hwl9/dwaWg6GNDOuvAb8fhZh2Ps8qAbZnaS4UXxBdo2Qfb4zr+nCtTnEfUUmNJEzpiopy
hmqCQA6efhHSC6IElBlrrKOxjb90RPnmcFwFo2m+Es3rCIfn8YSMuAIkZLtl9WRl6d4cJqlX6ozR
+ddZmnZZe0VJQv1ItcviSRMnV0iZnhVw9dc01fBnMFuxsw6jZaux9Saw5plURN5zRUYqTRplYiUy
5Cyo6bBA8jgEUzQPqeHVx+lo4B+BFcv788Qkd7N/IZ/j1KUNHJ0KCtTmGVWb9brbUVe/5xj/ugOA
/iucf5Egh/sq3dDmob8nKhsrmcUFJlu1T4L5kvQ5Q1m3yge+bUCEcJFOOMD8tKMCwbuFGnQhBATC
/aJQGtkXKeKb2LlThKeuKV7xxoTsAIMl5tP3Q5xFG2RW03hiJXyyqXJN4tibas53ya9dQ14o3Hii
gaZA+GVh0Fmz1qMnTHdCRHIXyo3dfiN/QUw3qmla3RTdOsYR/qybet09145BrPuHSSo5REJyho4v
PIKi2HIXC0XJWkdh3o++/7CbX3UB48m9kAgzbf+C5pDMXo5mtUfTuQp83S4lB0ipustXN7H26cPN
HwQSdWJ0kYI/9q8qBu/Hi8rcx2s3k6HLdUCAvVEnC6M4gAR/aMmw+yEPzHKolMWFYG3OWXLq74pK
BLMzqElocsbjQKnllqdDTpoKm00N8TwWM5KYyTROdancKgCyZ2a1KpnRwMJwS4DO7790zq5d1Laz
bCEXoXpnQB81RDWNQbElMujY64uHEum84KCl7+JqRprAz/KZXno6vAeUOhPPVeUF5k+YCHwmdHjL
5Mgp58zdtQRyfBh1KY4SAt86/8VupGDAuamHRYFYQymdb3/oxxrfSUEgWWXkkQjWUuAvbOJ9JxLo
zX27stLp1AsfAoPLQBhUkldt9rDFhKvSNkNgVo964m4TZVWQI0sCe/8VEqZEXnwzZUX+TK5dECLA
y0Va4TdvVBwYlk45tFcRHooImeJml7qYOeEES8IpFW4ad0x/QL8ttHyHWFJ6x7HDFXDxHX6vVW4+
VMpVNg860bfxCYh4O+872IJsTxRSH2oO58bUIytqcAgcruCXfvq4AgnHgOsr8q+WpTJ/HLxGehbB
fl5A17bIGx2GrjtOV96zMApSxERmLXF/EI7+Uq0oQGEIEqOTjKqKUZsPZqX8+QwNSi6EerEySJbR
N5UQK4PdidFrLkfpFue/Jnjjd8JbEh0hQ605cr2luvk3cWj/0Wpat883cKyl+jCrDtelQkstl+5D
FvOGQyr4o2JFDLN4VbN2c71lI7KjbAcCHrJguKEXAnRDewChS4SwjkgI7xKIbq+RXXEtoXFM9sOI
z0IVQyAxIGYFeMfGG3RbaseqAvwuBLiw1SIgjiWAlxrhoGkaswds3K9ueMGbGENPlV7STD0kl3BT
DT3ULwnLoAenQkDkrGWPNjZ85c3ZLzpy3aRkppyFYCSc6pkv8uvj8dHgGHQrkaE8A5L71ZkYNZeE
QZUUxlkZ4sBaRju33i9MicKh+3SJzP+jMDkB44c1eCJTa3T/mwdUD3Ga3SRz9yjbn4/XFAn1vtyW
noSZt24COS6sUet0Aza+mhk7rQh8u+ATSwrW/B6bWpY4ocQ8KZu87xX9gcwq7u3K9sK3Lcxwml4i
5OsZd2MUm1Pe5JOdeUhKchvE/l2OymYY+FbuNH8v1c2vfO95aFd5bFr1Z+HLkmlOzrPwK/3XQiVR
qqmidDdbondb6xq967rUEjTur0bPf3/ykFfpYAxOnalVAiH/H6NRxCPMZpqPolAp5rgYgkopd2KF
GqTSBq2ZBZHwUdLl8zVBstqHPMffRrGStrR9o8tCMNV1ywm6PbPFsA7s6td0evIdyHAel+ab8gxm
INQ4KU7RZBt8cKS+Lw17K1Qr7DkT6gk9xcupUnACnuqiEyUA2e9sSd4hJDvRjQTsShihCpoffjBa
c0FvcWVOH9trsj4G2pe7P3EXVOz5bQU8MZSh3BWxTebLVXDJ9S4ucBlc6oPhC/oVyazVgIdqVnLb
wS4CbIqjZ5O29Ltr+wuajcPRlKa5nw/ONCIWRM8GDPSNt+1gw/Wx+Lz1QJfaX7v49Gxu2IG1ATUa
HlSiOyhuLKj4XE3O3hz1/7m3WrvajKqveZisLFpvcCTdLB/dUOQENYEqlnlq6LX3gNqpmCn2UDpo
ylAsxptqkJsN+65hKnPgry5dIQwlSkNXrRkzAEJGR+sc58BCIlmsLtgorjXeyB8U04k8nb46617P
HNuispoVcQoxGzr97r9bhES+YKdYKs1UzZqvJpD+ifwZcBy5uDZK3n0BkNFrhfaOcpcs4uE/+R5F
KUqXDsRXDT/vGprjrC0NcjgzLwGoRF7B4bqo/xNfNjZwQsDg5rhhPW3HwDaI+/HGicgn/3ZPUf09
2qeq1BrFTEZ8cUda/LV2X7Bcy5EWlGrFnDScqz9JEkfltxC0Rcic6o9C9n0pcgKR/hrR8/AOJXxF
Xw1tODyGMGBF+xlffDFHZUbQpMMoiibEJXLbsU7RFZXie8DRsVk5u9QFndf16RzRPDVPnA8nLrxs
yPt5h1HXKMFFIODRwESphvvErwpvQLtMMW+a8+o+BMnGyjDJoiXmincGD107C0q0KxS/9tK+pxmC
UZ+9u2G69Ir11ETxzcbRWl1XE0Itug+6omqZsBKoYsB5jr5slpDm/gR6ZU5CP1VXrTjr4OIiiBpU
EsPPnBE1q2tKK5KM7WCDdd0D6ExEvhZnMSxFVv7BOCeI0pLW2ecgGOcj31Tu17xapN1o7LkQmu6h
U8Byuzlpr5nq59vKgpVYrZMj5FcJkF2v00QeNvmhkAiQ6lrrttJokUVUcuvbcE0tQZ7pFvA9KLSh
sALWmmgxDGzzN9psG4FUqUiqLeswHJrCHVt4rY8u/wUfk3fV+ct8HArk3jyb4z2Ev0n/xwWX4TXF
Py6E93mElsfSL4bbSN/zA+vwsqt/ox8RiYaeU9qt9nGfdslvJMpoBmmYHgGX0QBwi5Hkr1uZVuQw
4x4fY+h76624sTNqt5RGYY216ZYjHlNvUzfhgvgfVcAU9JAS7fFuGGGtpXpHBJdhKddj/EASNEBZ
jLHmXMJfey7WkHuyJMoVG20toq9Nr/tGdugAC8N9MoTVzxXlTUREioQz0dfC9xwwLFQ/6uhcVlnz
qLsPpDYGJFy4bGFwcQxivOjYbHjuSxERQ0njb/M/99Ql25quCMVpzd4QjzxFYkiXHHhpigQwfHsl
irjPSTd3vUYmpcl1aNj4Qmti0xE/MznarqIpUZswJ3tTUZg62hCoHhbaNJjnxV4CALKCyJFax/H/
SRdrdQGS4b7jWDPWyXy6Nm21V5/XxdSeoeQhtF9DphBoHtPDSqR4xaCMuwT6BH4CMFMRtSJC1bLJ
JnRX2cH9w5H0dEFG7+atjsmbgZA3JDMN3TBq/PsNAFIdY9Rf4IWpZhl6wp+FTv8bwr9WjvE/srsP
bWpgNSSHAWHnZqgvA4uhPXDmOvY2gnYZuWiSJH7uQxQtHggfTrUlyixfYEXwB1BGSLIPn4PV5Px1
eVTTZ5NkMPh5pOo2Y8RbhaqB27acTYsTnXXbi1lYJNYBWJamFMhLeqxRG23RwkD+w3B71q15Gns+
a5LhBCBKmxhJ7DH/Hb3fQJHQQM0y43pc6LZCoQL0Ut/5UvMdwu7ckAbxOFaR8nDJ/8qRCOY1ZHr1
jwR+3NaWx+Qjlcx1KNhXCyFmdXgWkRHx49eXIjtH7Rgfw8dG3zO2r6DxV36qcf8r69SKrfpvZ25l
PFg203qh42qFhWpykigrS0DRfPC4M0Mku/DbX157vFkUOoZcOJ5vzfcghgv5p/FgMpfej1aTKEWn
HdiSCW7smMSgOGeEQek/65H+1jhYZBiHYvASdcKEyidr4qkO35MtMWiW5yppqVsyiF2Bv4jeduVZ
F7G3LQ6zgnkY7wEG+G6e62H7DxpC2e1aeZrqHDk8v/X1KqCT7TeJvlj+38nldDbxq1jFEIXth5B9
PMoJV4mhKa9TjlUVLo7uchNAAdYKI5RA+w1kJhYsNvzpN52Td6PR1Ei1Vi1nv899GFnSWaYNv9Ii
FgJknXU7k63gacaVDkwNQ+VSclkT+yvfwJj5neOIFfQLxXr3q6r4KlL5zKtU4PaZqZoASZCF2fM/
A4VbMVrr/IJntpABPERlag0x8UwX3iDhQvAC1QViRVlbF6C+Qit3a+MTUaubUYg46zSPUbo0Cs0T
jykBey/VkVDVMkGTbj0rm5kmmwLlTC1lvHQCwdKQD18w+odFiZL2CkIS3T9SSbJTBz13vzZYC4cD
3u9a2MScQqrH6+JJHXGQgdb3Yq+paAtQPOkLSbEZ9H1zVB1+ygHcPISsCJXqtj7mXVK/QDFzI2UU
zwzuhZbPIuFR4UG465WuxCJJa4WP5hO4wR4jlF2ZxbrsyVVcQJldP8iW90sN3j3F4pjj87XXEkN/
1t7o/C+lG2ygOYYpXgkWTvnTEJw8ZjazeQLbpLKjBYj5QXkw9mNKLSwMPwNAkZWPvytkzrD0NAuW
iA5XeEr47hZDrZA3Zia1IvLKEpD1Zn4AomhO6xW/lGyzTKWeqBAITftpB/Pi6eM8UwOkC81SknGv
ANlGVwoR2VNUM0qTgRAa6KtgR8jyBCmimEZH8k4ONYV3mgFrW3a8rliY3tetoA/cqJ1ArFEWPO7N
YQExFhvkwZQInyG/W8g54hYbmJ36wHHGccCV8OpyXQnjKQsyKDR9YOU5KudrPiprvCApUEi79GFc
bXMkuOZ40tP36tEtmn9EiWl1ssBoUACFaQ5nAElwWKIzNB1zwWLuo8C7SKD0tgrRZiMGKf4kma/g
DZt0nWBpqg/2qf+dM8ECC7qJAG1uKrxGPed7hTaNj3og2pD2/5UtoW20kFJf/AjYUFz+5/241kau
BK9F47U8Ie12LfWDi1nvi71yEX3KeDxxCIIEtnwrC6yHPULB3vuut2xsiigUZmyv5H8iDOwJDmYH
ivp1Go7eEDNLsrFp2ENiTLo5J5PmU2R300C9nxtEbgPE7LGKEkRaGlj/q9nVY/tLKHAe7lnUhk9e
BfxFNty3HM40UKeIeBc4xcokvmtw9tTJtN1sMzMreQ/mxeLy2CGHaBl6V0rwZv/QFE8d6s3IMAXu
6f9V0VMrZ6JeKKlBc6nKxZ7Pvgw/gEBfPl0vOWxMmTpJOCNWigVS7ZVCB6f0pteK+scnH+gFT3SU
4mVv2Is0gWRT+3+ZvFfoPLUAyvCdoOznLA6SBupPL/Xygrl09HfLzFlZe6KMTchW+fcu+966znax
GuQ6I3nYb1V0FBzOr9U+zZLoWmllr6wa0BJeXS9KCZem6je/IcO6EgLc8H4uqYAy4TYVf4u1h57c
RTX0KMp/o/bESQO3GgeMh/iCJEdRZezIVqPkS6/S2b6SzJxx56Nf7BAjOeeeeta6gHJZoAr2n24H
dgjGf53uzppzi5xfBCPulcFO08zYa3bap9p6K4Sp00AQSfxIia8QHdqJmsx/mlCdH35Md/kH4S/n
t9ECWvd1WZ4BovGMqXyjaYRJ69VpJD91eEiDecPVM7kOKNDd9gft+BcpMOFAo6owXZ//w9R9pL1r
5Kd/ITkejhGyYiYZUfH1CA/DhKOmKRkvLeNObYvyMdskt5yIlW1p9iO1uLFKy23Y/gsnaXzK7QW7
gWLYaEHyAr11i1kKLT3iZEeEa878358QoSE0+pmBrDbkK6NwC1VZKJB94XbA4FyanBWmdcBcXahz
WLFHm0L63tAeY/MiEGiGgo8M4qU8S1vhaC057Nv3xoJIL7jwlwBesuTurGdyHoQfAQBxWAmK3MT9
rmIG4d5qVHCCl2cPiiCeHNkzV5qHPfwXU/lCC9EPfaDI4s2Rm++xZTjNLU8Tq8YuDwuRoA4UTQQ9
tFpaT6MwSODNoxVTd/h+vwd4NQFmTOXOkwBQWppHC/QzrpodZmeYTX+ZMg5X3ud1/pMWV2b1CYHU
LVaLTH/6mMxzvrX4iamrdLZfdedtp1sQ2J/9twtnIByj7wEti36dp1IHdBKO6v75z+wItbxYrB98
stqPTJzhK39XKpumzjgsR5oUfONVaauVwspC5YJcsLEtWHaLSz84F++chNxxdwZE1gvps2DJZNoa
EGE53QxiPcxRwSu+U7nvIy+lxSc2acHDX1VReswOEXHxXsq1RHGl8MuH+aWqEoqOdWsCp3DdZo4k
C8HDQAOfmeSH/AZpfbrX4JPu3gDvo/899iyXRNDI3LTGClt8PBTRw0m4V4Rp1uEWcLX2lXmh4QaE
ASduJojlQXcn7It7ivj5SVxsCHwnaRb5nGJRFmYjNR613ERc3xxnHf15McGLVLGHR48638oA/mRj
jdjXs0lYoiJ/UI+C1P1DJcNK7mcQvRSx0wufc+qx6CkLwfnNvUf4DZDEyc8KRCGoKxyjDzfjAzvc
WJlUnGlOq3Fm3xQZL+gtkZUiU0ZDfzmn3kszR6C87z7TC42Qad2wPwAG4/77vk8Jt+BzeLQgprYl
hVffme362/uLxAtSuIPBHFad0a0EElTazv4Xat7GP53aMCwiJG9M1LNbk/K6slWH7S+vIoJO1+K8
EUaEHdgdXZKhjLhXKKh3tXesksO8ePzwHsuTPs/ESlyyP8E0WHdnHDRfarTKm6+kzIqJ4ak9iZ3b
02IpBipWBOlTqOUJAtE7nijPkYsa4+mkvcInL0WfLLbh0SgjhyapU9bVwRWY0yrAqn+BjBQuWuxd
Z2lMILhkgCTQmKbPZYWB87GC6onCJOqAI0XuGEbV1dJbGbvBtEXPhZ5HFOxknLkhpmNUm2VxIH4f
I4HNRDy46jA2XZJWFGTcdpNIrOakqqEZ6yQ78zBp0X5JWhGKdG/Wdhsj3LUgbcEoLsErVLFVYCyI
+ijGmWBpC1MNYnVmuty7hd/wiU4MxYKnWDxaQfdOqGs7yXq4+/t/uH1qIgywRkegt23uvoffZYz6
X6j66bdvA7lj6V7FWNrerbPodKguPccuPXNKzw/3iP8O21x63TtFH5TCRexgi7V54/045j4ER6b1
mHw22yOFL4VWHXKv/cnj9DyeYwI14ZkI0KsWcpq+Us63W5l/zz67FV8/jrTqK0pshQ+wRJ9LvnT6
t1cIH2mtBlriNNF4EOjgVncbKbMUzo9Nu6kGw5NBSLrMTW4YgAS7+EI+6Rf+VM/znASDxKU+m4ew
bSkWXP4ewAQvHc4Yll7AhvnsaQ3tQXCJgoQ6NZtGaxvuCmik8HKgPvjFt10p6jdL8oKUQKHrQJAb
8VxJTNTQTP0f3SxMxPkjEal6ApPKnHLsKR+Y6Qh+7ZtyJPFParJ5KBPk20JReS1YcqWApn4emLeo
GOyNvaREDlN3IGaDm5UQ50/mIeqENEoYHyXuww0B/SSF9WMIbzbbUE3FVzSfmTa+Ay9db0J0XanP
ViuLpnVY+TMEg9aTVEjjUjylbU8igioKtYO9Pt6Rk2z18g/3ZxJNsBGDOltOQOfOB4XnOhkdywWR
m/B7iy5S17+c9na67u1DjxrDr7OC8dsbG4rCfuLHUinurcD5W/MKucqGe7f/2DbS/IBBcm1wdayV
uO+1/gxXUKuZu0B2gOIjUD4RnFlwDAn8zIPK4KR1cz/eidf/fO7kc24bxzfreLpI2nDTj771uVT0
mwtuSqNLwiTEhkvCAAA/aZ8rlioGh7jAVfgheKPHl9aP8BIW2ozztBm46l/4gWdoc7NouKyKxw50
oD1m4nnGFB3ciGSy+23EiWOukggcQB6fuNd9TFwZ1KuRDpD4ecysTbVqujbTo9nFBKZd8unkAT/2
WpD+bT8QvzFM+g/o8HsON0M3W5L9k54HlY3QXqO4mLbutyCjHTeRPXEACHjZi6rE4t7EXfLyG8Sx
FMOQ8XNqw2gLrZlDqMAgj9pExGnvWeVuow7c/xSjIbU5C6GFM7p90CbVhOl1c1uqfdqtgP5ZxZzL
QbuybrZHhxTXmxDZCd2bn6QKzej0r+1mvGQXVrAU0yxhaPTBTQtjnwTjg7NVpNH96/R1e1uVz+Zx
hDvz+B0h2Dyf+Os5w+Nrguz50v8Mp2YeZIbzVh7uQ2pGVSnhKvk1BVSVMM0oCJSf3+Jw26l1aW0a
uJ7jqmbtSQSMnn7qiC6FNKE6oc4MN5uVcN7V0XMNFzjB8+I7HhfJK/+ckc+gb7h9VLC3ibvziMfF
n2yA8r5fCe/3pQMKPfY0CI1bqEeNhHErgGfpiQKjV36RsfHs9Qp4DeGQFtFZO4uRekLZ1d2Yj6oo
HAVhSAYXzN7m389Az1iGYfve4n6TjEVo39Xb5VGwpFLmUczsTCZuUz0K4xGSCT904PKWRZJW8QD8
/vozYiKammPBiNmhnpvEOvMgdk1zJT/lc4hUKsOKOwhDKi+rr13JRf9d2Z283tsHwWLeLUKOKaXy
egrpXa5GaEayYEsiGihKKE5mlx9QyJ2cuHcTjNmkj2XdVU2YtQvzrsQWFdG2xk4Iq0vItKkoD+qX
1gJ9GtTto7pn8XgMYq4V0XDfrzIy0bYQGeSul3lxoODCmEWi39YTf8DtcJfVTvZsZ5Fe8ClbYp2i
YsyO7/63IT9mK0HjIPWg99+esgnnxGVj+NiJuIlMlzJCEY5OSVdjBDthvi9g9QyLCZhfClApHeCx
HT4v+4Qu+Ol/w5ccJqz2PvaZggo7YH/J19mFmWXbUzJ8bOLWRtV9vhmstOkx0EY2mtURzNiK9jYi
/kxo1l6UzIC0a0sFPjrzjk0YdJVkg2LqvDtVWyD/35bCUW4wXaArUgb6C6R2LXo/88iPzj+1CBvP
8ACKz+qY7Zc7O59LJwABM9owUo+52YxiaQjhs/3KnYBxSigeaBcj9iFh7M4F/g2UShRbg35hSB91
WLpnhTDnMHsed0ElHde6gBk0dnP4GYTKq2esl6J6/pksV5IxoH8hEVaNUh5J9KSaHUNBUi4AcgPg
zYAjMDayuDxMEJED4k1+X314BUFaXQY502mEJQlaH8fcNfN1v5UsNz908C0jKiWrdK01+WF3PY8K
JpStJKRkAxMFqTV0JHdz9sNez9p6bEZcQ2/sFOj4ioQtCinfadWyhiVVsYWMDfeGMc1OL2gYH2Uf
sUF7MaWBle2UXq6CGdKRVN5XaJupdUmkUOM7m4GhNHwkvwQgBi8QOfKq574Oe+qqKZ5qaQrCJnop
fx2XOe704RtBohTFSNJxyx6LLXUgTF3HP4+IpR0VHTkSYrYqr7VZ6L8M5Y3mTuxwVzRkVoqFajAv
wzzQAovSfjo8C5AkUxD8fYB1cuDPFQyIUPybxr7wqnv1DZdMJVMq7P1P4ZPR58X3mVhn+aeUSe7n
d4Xgu8oumCHNRuuOWDKnYmtl4hz5lXixcUI0CNKyZL+zdOnFqzKy+nBPKRjFomyfYlQE3i6UQc0d
GrXfYev3GTZTfHl70EykzALOolzTq6n+isAtCOCOArEj6/OUuWRuGjt03jh+asyfKdwp/C/CVQtQ
kZ0Z6d36lZNz5W0VP5vpIlsU3BlHgTz+6h+yqIOkZARbbUZ4BfwAUVxFgr16tU4e+H25pW82vUul
zP0NwLfV2SSeKX3LCbDXMGsGNkLf3j5O4A1Ye08yOxQqJTgUCjCVRImCSMAM1+hF7KFO8seczH4X
5P4R2ZR9W/y0tQpcetlkYgbxoiz6ilR+4nLl1hnXy7nPM3GqTln5E/Kz+PoPC+FG9852LqdGfnH9
s8/FGDYJ6Iqf2/NiYmRApzzA385B1VCLtdOyrpq5lNueH7/bgWnT90dCP52RtYlhQYnDoV9914Ug
BlCXrCvWWipc+WgpSRPEw3C0Ve7QEZdkYuVQVNhH7LfPhcLJqcfQcPvAEV2ogqq2FxcZpo1aiLQ+
lfu94Z1R5NS6arS3D4s0IZngFQRSfedb6+9QTT5bQQD1nkBLMmrI0anXYRXqofwvDVNuZsecCYWW
8THhaerz6erfgyKwwbdGKxosXm53yq75Jz7p4fgXqejE6sKY/Pi8+ynMD9zE11xQFXdM3I0uH7AF
9ciVQYcGcOjzilXsjbL8ooKSProbE7hexbTjog2n4FHALpFNvcc014I0+pkub+liInxppCaD9Ejp
M8hlf5NuWus1eZdY6TqNZQ+Kh6PXEwKEISzaB7RUXhyW52ERIyux3Rk5lU4Iiabpmg76sFdAmmrx
bqQ4w1k+As1+ZOVb82BWO2RTJ6jFoBkB76UO+/Y5UJlO6Db88sPPw1gxzSykzJeq3t6WeDy41FGn
ExSf8MkwDsYcn7fRKvno9HIXi46OlLJmwOhxKNsdQmKqC6qp8oylkYJOV2C4YTQ0JOCxvIZOsOHL
jYWEMfUKYDVWeDrvLpuCczkQp4KZy4bgYTQTbhH3wpOORQj3hvdk+wtJoeC8R0TM6PCL8wNeC9cr
qtj5boL+9pOEM+GDXROnDXriYPoPe+y4M8gTPba3OyUF57ACrQcfdmdVgHX2ad1oV7RfCK2pG9Er
ttXBdR+/2TvHFNpqhuw60f+6F+NkI2OD7U0gLgkb4owgN9NWi++9Eosrm5vNB9S6QKuSqRsm/t3i
2ZE8qjusToPguXrNFeVTYb+sv5hJgF1A9OrGkc+BOhxTFTM29cG7BI4wu7AvV9Wz+ia/Cjoa50H8
DA4PgEjcio8d56LL5gr1+lqG4mU5gN6N1iIxhB3D2mMWC9BcNI8WPYmZMglsBoaneQO8re8TFjdg
t/ju8K8VWeyiYlKTn8FBxPbIMeI50JjaI6nVGJWAgVeT7FtJvcDPyc7vuIHbK5KZiymbshw0heNM
utCg4K1p2ZabeXu7JmbEyQ6QzLmDV7F1kmmWnh0vP3Y9iUWPIUS837ggtgwe3tYt9Ai+gCXkeFxO
rE3Nyg1qIsVZWKDNusmoD2yAFMoHo/BWrCEKwmhzAA6fm2/HCYv4QpXo8Z0O5EU8FrNB30vT5KFb
N2SuGWkavLfFzNbZS+ZOj3OeTXxoUsukE4PNmosIpv68dnTJH8auYmRuHtMQQRcLQrb3z9y2vDRa
mF1n+nK1idoSc371VnNIurkJmQwIEfmmx/+kxqTwaahT6VFoJxXkEnVU/YIuQv44ZGdmPilAt5lB
S7dA3c3hwxZqr+RNJgGRKAygKpk7i8GX6wP5kXBb6wkjjj1QjrrTAalWAH5KNyaV3JUez1Gr5quc
6R57HMfo5fPZB8NhSzLysyHmy3a3mR5QLE38mjTz6iQbLRdSApeQFIZ68oc+RdF3P+LsJeZXgPNL
zqWhu5LKXXr9YD+WHVJeZrct553Le2UhtRbVeQeTP+kobqLSNM0WRePeQIJWMTzJJsHlvYf7mv5d
g1bChkqJ9uyE29PZ2DUqLSeaJrTHldhWil87DgvJmqrhh+PppRRg/CAUSvL2PzpodWwtsBT15DPA
IAtiMl+twIfZ8bpZi6brr2JiqYFQBYxvUZiZ2IutAEVqf3cQbgedTKKHrPYqDgzL8za2ABgTkcjz
wBzQtPQMuvPIV+Hhs5ZFwsiuGfg7E6tRTushJou5If4V2b3CqVQFZPMeRZU1sMJCBA9BomucPspf
P1E5BtKcDZFPhrf31gw2RfecAzxRgYyRyYPK+vWWtiZrf1wezQpIna8KYgAf89j86Vlwy990GXHE
xu+LtilLWQNEWvGx00QZYlQbK55op84cuubKL451/nY15ewYonzMGUTS4l2iSBLdZCw+JCa7718z
pKYwsS5DOqONosIpi7kx6AIAVfDVMTjPfbMBMdUTMNjxxI+ZiHdqIrCyuLB9e3yMUqxNN7gVZfDt
gsUaI0lN9H7T1iSN+l4SgjRrQyHYN1RO0a2UIJJSoTHyKMplchHr/dBuR6cJFJbCsAyIpyOo+hnp
rYj3QmcABQf4E9+b4q2orm2entC0mtWwI2denwuXUCzaaxfF6Owg1TRAdXJiGgTS64mX5yJlcxGX
DF19oyiJT/6VAmiyXdzpBpW56vzCagomnnEA5QnQ4WegandMWYMlC+0/7dYf/JbbKzcYE8A/6Jhb
3Hk8cwJnjTYfAMcT7B5LI9kO0yqNd8SCLZGKTdVGbmSzrrslGeDzZWnPoGMkrvtZoRuCVb9erfrI
doCRpKO3DG1LAKKRDYW9scFOkl2OM6vljMV6WH986DcXP713cJA/K6ITaBMZHXttd3XHsgtqPvle
Pxj84s/0CxAz0lhRNMFC0WDC/qaCdu9rRKHQLFsy8rFuizn/wuEDVti/F8DojSs/v+0Rjh9BMevn
zdqSMZqZ9nfhVPkR3AuiHWtklycv4ImWQ8J2S7SGHzvA1PK3SuMexGuP5AaC21gM2iUEeWi+efof
+K50Xg2Bp72PxdzI5PRsy8cc9S/9+VxGz68u7u6i9xcp7ZY5JXU+PReSifr7xycwBhm2OYkDpndQ
1BmEeit1DC0j2YC+n246gbhm773Wt6RlIM2LtEbCeM2MpRr8WqIIzbwXVZi9JLrHaplNG0vHYD78
Jxt5mrRCOzmws3l6IIB11GVSx5z0nq/1/lq4EV43T0Y5bNMwRWU6vA5p+d43ds/VGTA9cfiBHMtw
Xr2NA1UrSK4rtpmIYjK3if2N0XI9nJxyjyxFWZlsN/q1mnA6vlwXN7ZPEHEaY+qADbOsk77W1PBa
jTklTR5LM4QCDn1PDt05C3d8MXo5TzFwJgQzE0+PA++TouUsbl4zOnTagVQGYbdUCAgOAG1oScuY
ZO78SFuqhW+F0mD3X+E9RQ6l6iFYhf57Dr+ARLyA0eWcuu83SLbUCA6g5MkiDQ2GQ1HzUFBK4bGb
CnAI6pA0CwESpO4Aa2TQXK8GxsxYq5krPgbac8ImMFes5dYkaoJu4OqlfL/iIJTun4wNwVo8UsXo
FdCuKGQ8sL7L75mBtEsShVuUB3w3WmigyYgcFiBeNeviQrYEoiMpXx33AdPmeIPIsFEgNj2daZJm
/oXOB0+IzpISZjGjeTl6Wai+jEfFgjBN/L4kszXyKtzo2l4U2DGgkhInKR3Kxj06FHVLv/20/QHl
XV7Sx5bRXcD7F9sEXJqWKftMmEPW68b5NSvKgHGUb/J9Hdg5tAKrS4uUClMH/XOsB92UUo5f9T2O
mwVDgGKGQ38olo7oJ0bbUDPQzzgTPtDEv9sYzyv5tg9BPoJKgT8GXJkIeM1cIvuoUZBlUWNw0nTP
SjVyGb084IlTWU8Dh7Mb8taObX3OT6x2VYDh0pP5GvSa4EtsDqX3sWorQnDu88htaNgDvLcxjx1v
TAjmoa7Mg6XY+E3aUhKp58vD3/Km7QK1eEmeA57E/WNF7IXo4r5kXBo8Ha8HLt/xk6V9w3JW7Ujm
hjsrAkg0Y8HsE3P0s+vf87GMkujyr3CvV/h5FepH4IDt/12cpQHZi1PNgAWyOjntXnQdDNxS+T+6
g8z2UXOliHlMFIZPsNBqRhGSpYSE71kbdvEM4pnFqPEc6NnJU+Z2Ft9kRfgfuq9VvjUja+v2wvSD
pkx6dQBrdTDMvk+eV59+ZHyhOic0ae+sJUtBHdYuX+wUkrp2WKyBv/wkQ7OJeUMMj4UwAgoPIRK/
9++Z2h55at8YCxt6xziws/OW/hGjFKc1ocsXmsw5is62kUE6TWrktKSvDeeMcCPAoN75Fxm4S+47
SWjXkpTXPSMLm1swiRntcRUo8S1cFA25wsez+wH6aKCzoFhN/SdllQjKZNMlasgSKGulWzVhrUXi
UImLxb7WkbJV5fQDc8WBAFOK4s90Kx29+NBMi65yWFbtQLlSs5u04CEM+UQBA+PAlSD9QILeUfbk
cU1X1S97Snr1T2WAtlyJHoZW01fkD6rE+zomfgPDpNDSxN2UOHu75L68pGybgtBOuccc88htDqsp
Now8z7xEjKb8YVQIqxciSssqgBB9EtPzp7sakplb+1uMhaGH88Rjd618okJRTdiLSnED9/X5rAvF
QUFPt4g71YmQv+Dv+/m1eVhRSkRkwNneWKpqIrG4gP+CdH+FxYbaUdJQhmmkO34ua1/rlAF9dOUL
NOFXx3Hme0kY9KGYolq5wQJRn35a01lcBi3weJ3RHGrr7oPhuimMuy+AnGyvSzPalF/jP2oLdqZ+
wzo7HY6Nqb60uFb4yL1VFRvBMqQ6HfTKLkS3NFDyL6ghGDkNL6cnsNb2eGSpXDAzrOwtrdnQ0ykl
U1fr+HjkHsvp3Ue25eQUH4KaN1paHoX4JKZC00+ELxW7xeUIHn5mkz0F2/PeAkKFvQMQrte3gGa5
JgkbS8WwhnVYASGQNt9Jh9TwCE/DhFP3StdOWJzrteWp7Eu4CQHPM6H5gBM0glz6jTTSpD89Awkg
2IWsqUC1H6kFnHQ4w0GeHPJMWLeh+oIAyIWp9XUAI+1e8bg8IZ9ieYUj6s7llafxmMxZk+KOQRlk
RZPLyOalzQOchkStc0FfZ80k2AIeW5xe1XvKQ7DSFCKQsaMbdKtj9FlX1I+eXlHdGv6t6p645sUm
agHQb84MXrIiOCeZLhjYRbAWEaR3K0zoYhgUYs2ClZ/MGRWTyNmjviyiflnukIKNfB9G2I754HIL
ePPLoo68h76qn1mGhzUv+3G6wsFStM1L83uBjMta4U6NdJSWiw6rGUKo17eXihdYQxxSaNRwPfVV
YFiEf2QoQQow4JoDLNt31d8jQA9W32AH2jnwsQ4zXMHRph9CkilDyR4nbHFCWXeczWmjuCkOK98o
FmXY1PWMfrKIuiIzmYb0xFG8tldAaSHVu3iLnGwC7wbm/BGggqunOvX8JsY1ihonv6bkTZ2ebJgW
R13stlVArxdEPdkEUj7F1PWxK9eAHKJNySVGbWydk5Zx6yoPsFiVkA8ozRtkcWhdSjGe/u2MRirk
tWyIhXrVmIwniN84a5jxSmHjypX6fun9LPvzc9IAi8kq7Xj9ySdiL6Zjyjrn/DuRyGigWTLXWsZB
bva4FHUX6G58MgPgfjd4DmDolyLtQxU/vyiYyBe7cgp5WCg+3h6uoTdFSh8BS8oku6/N3XaNflLD
OT7y94MwQF3CUJrc5cDWsid/v5Kew42n2OBcDa3AEVg9C7d2+OxYrnJEz1Kum2z/HceJH8ZmSin8
AjkaOeBvVtulKRg7Jbtf4uPzlz5bVhWmhn95P1wwWM/LpPkx3cDQ4RAFOQ80NLThxwYd7gmwwIOj
CIhO08kMDevtyHpKjcTqOx/XXySeZisKS5JyL/YA5c8zzsGwLE2fL+v0Z+r6gdi48wP5RyG4zzB8
tnAGQxvBB+vo9FUg4d7+FuTEDX9Hx9pIgDJDhNLondVFEcY9Vs45PK+pf39eoNQMpLlyCQ4RFrTC
Ldc6R1zjY9tWCtoX9oJ7S+c7uTtiMv2yw9HlAdOZy1DijC965wmsKSBwcPqMmya0q60I4CXJ0hQs
mkbvGFzqd9u0xjG0njLXajjB/n52kjLAlO1orTIG+Ukr7FqjBAJyaZO+1Ust7A2cTRBn4zY87jVz
qFDC0rosKkawwBh39PI4bZkf+p4fIYJBWXMOdeUpbIs8PUyDKrOXfwJ1bwjWNkaL8bDl5iCjG/Up
aXL7b7AVgpKBW9dP7APIw/u1izHmBRjlOd9UVfK5Yl3W5IgNHDZeXUjbR1+68Lzg2amSZVH8NPP4
p2YQTufSOT0oZH+URQfnIlfI//XtCtS2FaahqP5+VfThIVw7HUFTVTTzf9/aNH4iDI7rZ+aWKWc/
MC5mnqlby5a308u6GnG9gjJOKzfexQwlSueLMsy8g5ikc7hG82Xyx4VYQi64A4oxsG7Yv9IQNogs
GBUkm3DNwR1IAdZNtXA/WA2BqukV555kJPlyp0+/xonKMRweYIG2+6Rc0OBgDtT8NFIVP993Na4s
ZchbOkpLLKXlmFx0D2Lk8vNO/JuzLDI8YC4zbvRIas+w83uEFQjKJPMnanzvQ07vVXDLOyEvhwdX
ANGOmVjZgW3tKflCYhtSdRrVkdgyCRtI+b7fT9KI6NXJ7tsGjK9AjYVepfm6kiODSVcsqsd1GWAn
U7gEtcmN8LFu5WPUjVxQA2lIr2ai2uvEvWyRyO9ayYuViAf08qqq4J5eJPZdOijAkffOLaanFxIR
diEhcKqATeLbkX2BIslHwWr5MJ3D/FepSlJ735YyOMexx6sjwf9ySJo6xHPP8B+IGDXaIOvYV7ev
T1gAyJ8DvT2tRlTyVARyIiI//AZhv6dPs5dGAkJ2uG2Pas28e9NE4iwEfokZorzG8ZZu91e3/5nZ
JxjkmftTBmWkZEOVvVFyoR/BueB44zIO8niTJVE4tMOK/cWBa0weN4S8xZE1wKMuhN51wsL3nmUm
J0SHRLOcYp9oJyI4LqkNdg7DXdjzMKKb7MbXDOtpwfYPf1dBjHP7psiiWsmeDRO9KTv/5C8fDFlG
vzA8TX9BPM7gwtqcoon9f4YbY2p1vYBG5ekNwpJEfkLTfl33ocGJvhb6uQXAwdxrTs2orWoDVcx5
Dze1z3AF00y07wnbJqTE4zbbRZbJU+Ttl5X0xQ1W1FqaSZyLGV1c1D5xDLzw++8/EMYa1NzHH3QQ
EmxIJ609rKBS5+r0mxZQ73Tql7XhtMRixp2F++bfchCOeMX/geaoh8Evp+ntsasOQqNOGn0Sn1wS
naoQbUHYFF0ZDaYL2Xwr95dQgPPPvDp5E1AN4iuCgK4gtBtqU4OSwc0rDLZ6efLeO0PDiPTLr9ZI
PJOxSIypj8y2ci3R8Bzmek2LYHaP/Kqdwe2Zyg7zwjCtoTjcMM/6JK39EZPvUYZzGXT1Tjc+xZSU
/XKvQu10sGy6ATth4xYqRvBqxiWuz5XwO6SPRloyrvt5nGEVJLOCbEZ1VugRy0qX/LokmjqctKXE
4FtPnu4MGtMxSK17pWqhdJjByGkUSlDnJPM2AXxLOyEWNgBcV+GwsZiw9F1NGCddsPBttIn4CO2B
2E+5V9n3Iw0xA4zXnJ/vKYMbzcLLId3iZ9c5veNrvchMQWCppe+zp+uHSBHI3XTpSCYwvjLmYPeV
DExyjo7yet4UOLAjP146WCJt0eRuINd7mzQf83vdm/tBRsEW6RrmTeUPY7+Yht8H9UCgDmvk0RSI
ByEVorZY0UM0yJoyEDs9UgbQ+zk/rzaAkoGL8FEWCTGaMlEeNk7fJtWUt6BRy9yvmbTHy3+Z4shA
1S1NSHYBAFxGXv4Navrz6I+0ERfq/9qScO1OcaKSTzm1QhLK9ws+9Bpn3v0ww65EIG5wwywnyFnb
oCbGfCokwPI5NSDAbEtpC9TXZgO7g17cdFV9iIqtAbXXe/eZa0MHZ8jPBYlb5NpIp873mjzKhUbd
qTYSz+1axF4Zy1nafG2wfSNGjaM7hP8jZVMQl4cERVQ0leqKnXYDZVJXFpWeUm07iAbYg86JXhvd
Kt9+kgHHepPolqAc7OTBBo0a1VdV+cjt2Xijd9jPpjBh1eVfHzoValkY4VHruWFEBZlYQulmpr6b
2dUYATVwHA3s83Zagp7NxYeuPeAObi37h6GBhkFffbvPtUByeVbAr4cuXysmz/SVeTuQXCwbson0
3GjReAO2sIWwE2sI3MSQoBO9PhRkml8vNnHYT2N2uCMjaw5mMXPX52BDpoiGi0XNUXh9jE9S+oL6
cD+v90qeTaIQ66s3VuOP2r6rwsZyVoGjGELXe6NMGpH8i8xOLp2p6fUo9G5epjV9BLgzd4I7DZWd
cw59Gp9479Il8HLJWr45pHpxN0HhMQYjeBDTebyRND+X0njEmrv2fpd+6UrM/KS7jlG9XcZJvCvx
jjy4CdwD9TSl6xJFU4IFKBMLKapqYaPSR/XCRu4LTdYVcUY1WLNhosrPDGblasXWuYnwvJHrVKgQ
/geXDHhfbRPl5R9YLiB6no+5Kog/zZWR+bvhYz5qRQyNaf22GuRo3y0xUuMu8Xa9zTZ9itqD0TkP
A+E8IgH5VZBBuB/bkjsFlIB5CNynXrJKcYy2qVTJqZfVevukVdUnxYN6XUuMnYdWnpYV6clIgn2p
FaWjceIF5KsFDRtpeuOYfeqB768B1QGBDyZyZxbUX+TPr1/NuqoabZ5CaOZKC1I7UwBUSHscXHKv
znUafdnDN5RVl8CGFjwbatUm9uV+zM8TNfZOPfD6wlyHqb4Tu2WOL3KwWYMxULleIXnsvTxlxhzO
hAl7G0JGk6//Fu4lIUD0R84VkHnHcu0iJ+Dr2C1JyIkVB17hww3E8s14ogfcLN2Hk6214wm2Ghxu
f/jJblZt5yh/YTWt6t20O1+Usjug0BuE5I4VpNDvemUz7fIVhHT+o0tggn/urGwA5j36/WnNuz5m
8NLjWt43buYA0y9Ef+52IpPDmtrOiWPpRil8QIVVfMCHaubPW7EIVuyaHHayAAAVroYD5DekOjQe
mA25ETVVEiysYEPu1lx3Kx7FLoT8BbU0d+ZwON/JTsgVAKWVW9YXRzQO6ga34lIRgJQA+RP8UHaW
fzu+Vp16mXdv+Uo2qRy2cSk30xHiBpyxwfmrCBXxWsJ4e9FZNhDpeI/hYgqSRGnuJ6RftPjauzWk
qshOrPJs+B3kU6kPWrLN1CtMw4pcP2rQots4ynb/QqLmCPcYMnZlgcqJtA0/RePe5MWV6ZIdL1rO
6WRbCLwkhBIA7LU3JdKy0XW84IcLoN/52I0CXcjeggTirwj0j0IMTTqGioahpKwS/uGE2oI3gEAc
BGOb2YSQiod5XYlNEE1x+g4gYvZ8tS2yc42HZlTvjXpFVBya0oEOIayrkczCGvJa9AVurYIUCuaR
rAn9YMLqYXXlcWUmgypuhfeTKOFsG4Wnc+rsBXPiJaY7e5mL6k3z+iVYpLAdjUHGee8BtnRXCRBF
A3RmuWM+cMju8tB3b++I6zlPwe0Lei7vi0kZ06D7cH6kc9rAapiW5f2U6PDFpOAHCXCe5IfKOw+d
fH3DOMuhktI+ZuvWYxWDsC/RfmfsEL0ubLzb8gbg41Oez0e08Tz/wq73Mf4ErGY5i6fB6hStghGs
mAE+InLqLd6QN5V0Plbp1e+2a8jIkd3FLyL4lxMHKf+XuT4PUsFnd2M12q/cBd98vS788CUpjrBS
eOf3g5sGV3NY2vsCae1vB1cMN+F/j6Szi+XijTCXq0cTX/fz0FwR5tKk5KaF+kgr/tI6CA8yQht5
19TNYUXaHG2PaXXrFFdurTmzDEUoDL8bPwsydPm07AGWmOpqzlbq/Lkgo9QmxJ9vrdGq2eLWELUV
VD8S52SMumza3rtkDtgsH7inKiKZMOp/5+CcOsWlhn3JzhcrCj1Y5N97TNAXvkhmkUXdHmJIlY58
HJur+/KAXmd/50t5v7iwjxxYVQNKEBKP6ghXDBsT+17qtbco/mTeyxrItxuWthXbXL7jucSWKgkV
fAbePYpFO3x8zCumgzEWA0yYLVoKtnSvLdPNbFmbZwKqnTXL8kcXJN5FA22mrYaKzaxjrHV3BVsx
3S5slasvBRch9rkvjITklVzIYX4AVPb782bHkiRJB7IE5yoiQx6jKDn0XgifqjLmfei8qCqTng1C
zHKJ4EQASkrXbyreVr6lGGm2/R59kuzl6i0+4W3mZHKvPoJIZznZrcvenCFTMS20IYM/IucaXhO2
ddkhhpQKcJaEqIapPwa6aqvU7QY/xBlN6OUiIkSBR8xs7h7J42YJvfuU+aIRb5Wm3HnhjW+qHeLo
1Zhk9Fw8Z/u0fMcf8waupGNDCDKZzA8xvOnsiIGuAAS5IqLm0pHgMIMGjlG+TWszAaW5O5R39AoD
JcD55mJlfbChoYI0+OI/S0yDBUyhitCosGIIN4/bcBIVhsFluQ1Y3vmvBYCFYJO01mZs5p3TXj2C
hjxAoUqVWBTjQlfZ0DTro7ozw4tq8xL0ZzUBb05nUOWCfMmEzNP31aVFXXS2ujnE7dP1vSFhezIE
YCBKv3I/Q2Bp2RPDn2uzCUgRW8fdmCqFu3tAzv46vT5joiCgXrpk2d1Hl4xz6HoQNetYH2cTtkYc
7+yp+pNEo2Zb7FB1JJj6h7UD65aPb2txJGrHTe55aOjGX0N2plN9dhXpl6Zsge1ZhRSh8/y/9zsg
Wp9YxMS14iPdgm8oHfcnWSY6rdNV/YONlTp0BQgl3vLrZfxsBVWJAiSbH+n+LS3zRP5xv5OYja2r
pv3JxLNVkuTgHweK3jZgkpVBS5pe7OewtV3o1CxoSGt2OO8LkOnry9gtDUzqGLHmCPi6QxwGuGyO
Rty2ms05seej3wVj5T33zO44vR0DOhSdnZZZW7UHIuOHx7hNIHOtAETq0So7rmbkRM4blz77TYL+
TFghty+cQV3S30f6Esl4pvYUPZKkq+ZPd14uudYD3lUbaIav65pBAqcqJSvY8tM3rzuHfdywnrC4
odBsgYdqMavsT5nHNiwXY8c1SvOCodmKHzIktwHS4BypMXEep0HILXQlDDxAEfIPtlp8t9NcX2H9
bNqEIIuPuBYM0ZaKwIkdaW51ipeq6DIrk+BKbKIZHxEvYJ6R8e1oWUpOeuOwKCJPx7Aoit8gz9N6
PDduX6D3+h1SlH/yjQdq+jPusIvtIQ1KbiaUksl9y15bF05MmmTuCId84fG4SmWkPt1NIpTrnfdi
1s9wX5QPGTU63et64iq+rHhMJSrjjuxj4jlyKbW3sUH+236e+QQBaMWikV9bCKJA/tF4lNzyQrm0
+sXoO4VL745SNLlmClYsTY3ywKH1N2ipEsVuDOsib70ug4IP/5sD1ma5YQSNOSwjKwAvwn1nyFz+
3vT7NX26PwfMeD/QpHgcseuBTWSechiesTMQIg1JJzNXlght0LKoMtAVskve/mShD9i3TY9om+l5
UJXs0DNXUsZWfbW2vmZOjdr/SJiJonUOLf9pdD1zIRlZt7U5loFUtRAmmpInWQauSalff3Z0Fp/u
3Pgs+HOk4PtNoNf3JuCsnFhVQXcCaA9NFSDcD8cWpwA5VlREly0nouUjPPdMsVjliLo1WIZN/ySK
6OfiW4i83ENQjmoYjUQnb8xlmZDMdBPONVDtMNlIHdsEaB7TQ6xb45RRbjRNwSjIyQOiQE10rZns
TmwLH/ZTO9HVsFec8YqlDU4yOC6LGgIU4+410cT02Ipp9szvikZUoR9zagYVij7gU704F+rd9If8
MKVnvEwVVrq0RpcHtJHTOLzJIcU+FUy2Cw+teDEIvRois7xQYrueS83J94c/Rb0zW745Toef4Ji7
XKo1llzXRVcf8JKYKzyFprYKIGzxIHOAudpugLZWrgd50qXnQKCaKmOHP/l83OU3iyJmVsqE5zV8
W5MwhVf8QTmTLm/yKu0H4Y49v4r1zM0eCXBk2/d2EqaAHA6MEA5/fiTxvlAV8bWAh9sFuUdlkzLo
9qcASrOyE1uRkBxBwDC/Yww96l6jN50ifI3x8iOyhYKG6oYGnia4Jy2RvF9X2wyOB0bDFPXxNCoC
iwcbXSyZXyz3R99wY9/CWs5Fimwa5VeX6GDEwDO4Ns74iHyok1YVcp5Y2kOcRKyHDhMaNHi9j0Sk
12o4vJaClDZsjygxVSZr8W9REUirnVk+pEWbRfhGD5Jh9AYOcHnXfUDIsqxLwu16kO712Fo1TqZ+
24hr7sdIpjo+aVmLu69GjqVVCyVjidd5QFqcskpFYYrkO0Z9jk75K4jGXS83nE5uj6UqMwBXc4T7
nJYmXdR8tSh4bfOTgLIlJLC6F9XGAzQLpt2miaQAaCKkjOvHDWRg5v2hHO6RSMDJ7lf1BXiiB8xK
GVnZZn2TGmYFbMVWD+7iQ9WS8La0eP5GJ9yaZiM2hAvOHX/YfammKUTEDOS7w9I7OYI1roZxcR/7
6zaRAVU9q4aADfpcgUliWYsj26exByoJBGEf7ACJWzS+X46jh6CRdA4eHiS+dIMrGkanoyBNvQQe
n5iuRgC2FOSfV4I4p4Y60/Dtygp58bMBmqd2sSbOQ6m127l4r0BPWa157wZ3OLP0Mj1A8Mz8Krn8
wITGVHSgzl8qR4568Bw+80v04Qz96jZjeh9u9uWt8R5/kvZIVfG6Rbeo2JeZpedLyrWgUXMuL9VI
KIOEfQdsrJrGB+IV5rJy8se8YpQps+zYB+KVMRvhAWkDeLePtGvEKngcr6ibmBsfcJvb/nwPOc+s
hjXkIuj+gRoi0Rr9zD+O4kPZz5x4eYI5ZfctVCWnnG+QAA/K5RXBXMrYLX4EZUJjl3LDhDfBsEhF
ZcezJUU1/uA4kihMpqxrHwNQ2DJgU87XlwUSNSQP62Pg+DPUP9CN3AF3noKYEu4jbd0fGwevkv/L
amPa/Me9VC3wF0E3lAWq0E9+0JJdUvPRuCGzMZNLmEL7sjz308I30/kEBHpCCE1rXJy6jqD7J4O5
TvHWkUM1a+MTkku6iZivDe5EKqZeKzuvkYM0lU8uh0yO9VzmxnZaahv9FgQp/cU48xzlQZ+Tayyc
0AB4+e3vB4El4Z4FXvtX4n+JPEU6YFfxIVAy4Bj7A9KsWnhdtCiBIBWnzM+G7KNsZwUf0FSeIEJM
2wov+6mWNQDD2VlAVkJRBFwl6X8HHXDA32JKpHcKl7a2X10HU0+pOLmk8EjiN19WT2wd7l8w1x3x
d64VE0Q//ptjI/YuOaAQqizS+JJnkljXd1XCPvlOuiqkXBb42OVQtgb2lDB4BgC77eVTSIraBwkX
67oO5/vtHioX6097mqht+74bvR+eGo/RVj1fOtIMvuWok8V/f6oyHP3fACBpLA5a8t4hndOECDbS
m6fvbTxJ7WkN50+NoH1A0OhkuZMrgl/FNMkg8v2L9LNaviG07T+X69Ve3AwApN+pAZsfyZO1bAUl
TIVQRNbyzC5zmzpG1UPUsUOFaquacvs+3zbp396dh8zlLXaRiF3NLCbFREzdg+Ebj0LUl/MkL6Yw
QWVMVb9UnDEIYFSWUNhp9tqBvz95DBXwpyBP6ueMXgb6f3ZiAU2H/9oFDM83dZn508uevMvoRlCb
atamgpy3oJnBSvzrBJIgK8h2StUpCgwgJ46mMhO3vxsSgh0RjIRdFpsCu+fSn/3Wxwym3bweAM/P
NiAcCJQxgPveQ2qgiH9hlZb1v37Iq0MnhCl7glRjCiYjegP+MFvOEK2Sm4RW9aOdCrezhNFRT5+C
DHWHoqdeRC4iAtiI3agV/AQOJYH3T37rc0d0n8pskoVamYSu/mvoRxEeO+qPoSVCrm6k87rQh+iE
G/AtO5KvGKI1dd7cSf0KyIjW67QeeFVuISzyD8vNC/ITVAm9XjPcRYnjtCsdZi23MHVWIka66r37
zPsUOZHm50EnKlywQpkeDzBJnItXkJin+Xln5rI4spThSHRtb1u3yePEFlT8yap1+bQhbOVnumVA
tEL8+/i9szJTHnjEFBdrVT6tBsDOwSzjOo3OeXAZTFHECtqEQYvn0E5Bw6gDSl6HdCISuZOd4/w9
xBiZ4fv4qhmKVXxvKiAuSBVNxmVuoV6Rwz50PCaRQtX5I7Mb9yzmF9Mb2rlQmNXt3XWKSfNxj8F9
CqwPLC/5tM1YIDVB2OOShro63N5Cj5Iq4d4HYCchA/NZw1IzXITWPT9w16QYt4wDbxn2uROWt3yU
G32Jbk0dF3/WPfVd3eDuhANby0saxZz8ZcTnvghcUWaaYpwHGumOlDQWDLm0l9iFg91UA5cG1dVz
zeL8XyVZfBv9M79F6g8V6KDi+pGeF9H4CPmFiHXe+4oHxFjbGSF0hztrROzOwT8WZzw/L4g/yAcj
4o3GCTS3lchNIUazmII9u5xxT//YNtpMrnIcYLj08UaC6zrJfNNTmZkt+zuyRgP3AlhKtkbbRwV/
YQlcfu77lGKOPcZMe0XEFQM02HdBhT6zO8utUmhNkf4OnYHSSJImKWjfw0Cy6UICDkf3U6tlGJqH
XcvYzm8wsGKMOdmUqT8zFMk2mkVpln12eI4+IbZx6j1+jyK+IDjOyorJWwrVn28Cg7EEeZuJRCKm
zAFTDnK3+fg8EB0NQho0js/AzHTLpvpqUedAE5ZzrvpZh6moxqZhgnwhYa/Y/Fxj9sr5lAL2lra6
n2fZYa7JvHFNsnsL/eLBb/k4uib6Fxjstj4RNXEn6F/aHmSuNhbe2uRGzvU8r/6gaSharbZvtE9u
8AlTLAR5lWtMiN8OeE5czipfoSRCtx60BmHJloBaS1/he230+l7fqW6JlVfMpghAT3vxHjQO1aoK
PgrU3ZVqZmUhMBrdvNzubLh3dJKuf1P+BNPNXVUueNobx73YF23UqDz6tfhpe0RbzyT+Qz4AAYp/
yFLw7ZtUYUwt8pUCLIAUlUIML3MyvJ7V6OllpkcmF9Fm3VTuqA+U11n92tx1LcEHFQj1Sf6g7mQe
PdQVf+zoYK3B+MlpKpUx0cd4J2F6a6oT5D6tHq0o61BwTKN8YLChNJ8tTPG6a1Kq3XVvoOgSa2J7
oDlcPGh3nC4n+edSlko+YZYi+mdaIDm4gDzvusfpUljXzdWYk8VUuFWnKzi3dxTIP1aEKmROWEfd
iCpS7PKE8HTRc0BiDzO2EAPgievikoI1amNhLCTo9+rS+GMapnL6NlCNhToUqCrT2qRrIvAMjxgp
WMUm5v4nDcqrrAO0p8JM/v7AWhf0Gz3sg3FmVfTLvsDgoaWzUVjFWdu2Q+niHEAfOWmyi8BLoSBP
kDhg9EV2BScr31Ed5QsmJXHt3+YSk0vuEsXGUwjBIvjiB3QuX2xbTkbVin3nYy0umYvTzCOL7IZQ
y3tRqmUIgLod/2VOVKh1zCqvrpZjBhnn4ieTWAtx40Y6wSJOQBYDk0i5YY9/EqBI+Flq2q6FA0rE
dUVkyxGHOWqmHrX5iEAlw6Esyjr/XacGHAsQqiwv6pY1nezy4ovbDQ70KOpw4exAAP2T4zxK7Lvd
V3uxN46XY0+zOVeVptVX4KvEuTj0qiqxLk9FlkReNa4YVqYHCk3HHSz01aC6KS9q3LMBKD8iyuXd
sBtB1bPbstQQF4FpYNnlF+RklhMK/wVXGoXElEpd3bmvhF8EQfuF9mDuRHnr82EUxbMAXcZeGg1D
LaGaEFWtXbTNtKsMBfHqZMgo/5pj/FDsVZxlBr8ZRRxxFB3A5g9bgAUQDr8FyfJRw6Ebhm+yCTBf
zn2utgn+vgUnfzEWoHEz7yAZcevT+iMAMwHGs0fWXUxAj8xQgkcgPqHMiuv2vzPZzm9jMjuXTMIT
+V9nyBXfQ/7EwcVBZBm3VTTe9IjCF++xNrNSFPJyd1vl3qP7UPG/wAXI5vnfecH8OBeLIGXV8FzU
SCt0rAIU0cPUZaTgWdOZRf/rquXDH7f06APzdr5sQ1nOm3kL+XMf2nWPBYubL0NNORXFQtXa+Fvy
WLwRt+SfYBeuy8x+ssqhO9G3ItUi/WVhRphR4rjDFOofoYXx1YjsYxNxbZAKAVSN/POg1khR7wMe
PDMDZtVVYfHoVnuvZsPMLNdiWcFU9HEtqf2d2igLqKboaluVGSy7/xHwKreWPce8gRbjF2Z6l0vr
Qbfu+S9JCWW7zogB2W3Uy85Z5k5X9z9tgzdxaVGcw+FqGA9tQuK+lDkAYkcc7nDwiead8DjTwPGT
fPYc2pz0M7gtnWS7CW38EaJjT1i/ilMayDULkeG/2zHwtTfDasC842iVdRcE1ldSbIyWRJCNvqDS
F517Xze+soVwIbBAlSsx002gdFDmjK746tufX8l01pCbIhBhLQjc1+0Rx1WOlABHZmB+HmAsZ9yf
LD8H9EQdN5rYvAEd2CxanjpmALnDRZhWOGlIHGzHfBDR27aW3txLRlUEZq/NUprhmAvq4A/LL2fC
z1m5YLmWMt69FyZAFFg0PHFsr0PWC1g9CDh4KklyOhJv7tYKLb+6Wjy53GkKt6v6TahqIlOxIDlT
tez0rSAVLJAGOemTSPfKhB7BqMlwQ1MIDkly0FhXeR+7tvqRv2sgT5VecRPkM5jvgRDhivExo1aH
f7mAMiXvan10GXLTgKwMmjJeAueBDX1AhLLMc+JaiF2ojeA0EE9udB0u3JNBB1n9rH1qp4Vi5dqT
zWMh9osyLLKiM/r7nAPQMymHsPRpDaDOcHZlYbo15ISecdEc/UCmdTR6yhxvEQRU1DnjjfwqHCpl
uwEWRpc++yUaOS95HBdoP64Q3UAllArkZr1p9YCmrhD23Lk8BPdWmccQAYrHJuwHrw23eEmoRSN+
BGGxFhMHBTS7zFgeFCdBEBm0l7fBZLuKVzrdZ/Wqwr/fGhNuDTo3jj7DxktDuX+qtHUKoTkiYzHl
V4IpsrCSUM5RkKZvuxN0MEQVaMrcSckZzSXIJLbYat2s0fSS2S8Hdee29Qn9irsqinRRmFn0CEIr
o+2hFI+d/I6ljw8XJQVg6WhSop7pQfLVf/RUzlzbM0yFo5Ghy//nr7XBSTYjLPjMNkBP8axNqJet
qGwdMa1/hZvXYpWH/Et/o9qC8cYXP1nJWqAO9AqePSFY+aoxVbFUtgD5NsFTkC0rjRtxXJc8sTZJ
ZRIEHHBo+IC2pfqBaUlrAWg3XHO9xPpMmFtjD2qsCLCM3EGFnG375RQpEG4FM9O4Un0wtIUuSTX9
TsRKe6xuPxfQFWp0QHSck/fs71uHkSVAcTSGHK5dhBD/EZb1oqdxCFGDJIw3dgEwfHRgNUW1Y0o6
+IFQ+7+g/J+dmedCMx8SMqgyGDTKqlHBHHILbyiVEeVA0untqfYIq59kfZ01Mlaa/IyexMrhVBuR
7WhydiiTr9eG09Rvr388dV8Dr5rnuXB3Eqm0W/d9MGrNTFnBJWjq9Pgy6+2y64Vaik7jv6WjaRW4
rS8Rtmd5PEGAq0mUi0JJTisK9Z75vgrL/l6MmYAVm67bFtOolNSaMCOw4XWbOllt4TGk87zoq0Q8
2skxi1i8uhAzb25vVkppxIZ+tPS2brbyhpgPmUnILMKfhUzyA58Cizc4yDNGPF2HpJwokUJlEb32
N7nKPvBb30rtwFg2EWgE6EAohcdAn79AI0tLnHddGLK7rvthueeqV8d+rPmYqUHT1ccntuzUDY8D
4StB2IDCj4wFHxggu+kDN21x5gdI1G+6flgt2Lb3t9CDspBPQTXTFZbW5mZpaWuPLIr6BtFe3gKX
dPnyqAUznAYppMYV79M9CvpWrEhsvlfnzVyJZ/Sm6bOs+hCnuTr4ybmsH3jkewxT1yS7n8lD5U2u
1wiUvocX6B1h3QkxmphMYA/gjBE4FAxX5Pzz+kvPl4mEcXs0EZY0wSNWLXusSBJ76RBd+1m4o2pm
tOfinPxQk6gDZat4heqnYAoLn1JMKewlUST/9ACZhenQ9CYeKaAtX1dugGBxIHGtrkaGiDRypTlr
5EJnbYcE8VL6iVfHx/QevoS3dZTFTOd+t48Z3YiZgYdu/0akR5YwgXdx9HfhWOt6IfOJQ3yvFOnL
typLIBKlRyZ9G0KXONZkgyZuw8IYMTVJ2Mv+GXDLPvsw/lIo0fFan5b8OcrHrz5pQ1vpOmMd1Drw
9cIl/dINq51O+w2LViLBT01mF0rey2cwk2Q9MOwcsTPZy9Obq0Te8VwOyIFnUfz/8VBzscoahfC4
uZGnJBv/LJGBIzIQTh1P2hsNvlPFSL/rmBvqr3RjplfewwANgQxI47ROTp5Q1glfdQz1s/Z1M4so
4QquNVKfV7nlW2ksdp3O2fnGnnT6AHHssgHJZNMg9opKFrEp6ONOrVIMc03b5yhkBtDSrpfPGGX0
MrnHyx32mFDbP09HE+k2Dc7asvJDhvupXX6mbckxfDrnKkD9N1TX2z4L1gemv+MYB8L/NuH+MjWZ
mpVUUji+QVBy7BG34cGMxk/dYbjA7UKQkLOh0ndMkKZik+B5hQvpXKFwRF8ZCaKHpgMr4cijw+2r
qKmrmEhnStSTzog3SE8arOr2rYvhItigVHuwTJ1M5KI9FxOhwZDOoUbmOv26qQr8AlS4e07suIUn
aHQEpmLG9p98LIHKdfOaGiftyM4L1mVu6hWHxMeiJ3KLEZK88AJGT5i0dESS6kNSkcTApQGuPu/l
kjj5LiBYMbB/O6jZUkC/ssuLXhQtbNHJa/R44PGLkehMzSctZawb822lkdWdfM5XNJNk6ATqEZm9
K0VAzRzWK+Jcq4tUiJ6GPmgytbgrrIkKsYnjCtSKXQEVaZRhEM3B9BaIEOLc0GyqW8iEVUoEc/MK
Y6eNCmWS3bZzYSAkAlBzbTmZuAFH4xP3J8Kr+ObKq2vu8gQBdCQsNXp9UBfzOMjaBizD7HcbLnYU
1tygfWDyCes5m87o08t4NWXau1jHY8TjrYhjuGqlB/TIoj7EIok51V9gcuEo37IrZH6qzRm7mPOf
3ylcTilLxWf3j9Ix0j+9TrgPTtnCJaMUGp5XVR0fxNiM+FuWmY+dZYGWJ7iUQtklWfH3BYSn6CfM
WHDf949hHBnDwiwgfR7RKP3blNQM2IerNnbN+FSGnbsjUqxSw7xkITl3pM0+QpndgZ506lPTtYH7
1VMlygwxxEVYHfKU1fh614zZ3iw7RTqq5IU2DO34uzkgZTchz/OGHNK1SA+j//AtBAl85WHktadr
rllIDKgJ7JqzM06n+1FjAlNMLT3Bnb3WaWK0kHsUEKVIiXlLwpRMAN5VJqpCErGremAAvtZ7sYlr
EEmWcDMF/OAj3F7sFxTknHPYSidCo1TMd2ttsBKi157YSWfMbTFYZf7j3i5+mYX7enVGQJW+dboJ
Czb6Wk0bvgQL8PAWVgQV3ApenLDlHASc8UKIRYtKM549eA4gXs3cGLbW4Avpx9wR7tNkvFQrgxUK
Mj8WTQPOTvjUHbtV0NgHps4eQNW1io0XEtSSIsJDL0XZW7aQvempjSWz0iuKUypSOlVq/GvA2MhR
2bwGIEq2ZV53SRf/HShHxBdG60WuEsIRA1oY/6a9kRcCgSDyN0LSnsCwvzy/uOi8AHQE1RNOXPot
gVrwsIGdsaBUizo3mU36mKg+Xd4hevG8djJ1y9oMVb4nIjON6KWLr50LwcJHvO/oMgzIfIM/srX1
vMh8zVIR9OYhnwYRzW6K63cpNDg2OiT/0XqhMPkNjpFuQa7Skg1ve+xbSCSexufFRniXcikzFZ1q
K4BpSPA4WHyZbAbmh8nS7DcYAMkncx7t07BUsPN8yS+JFXqvnEPOsHSmpQUBCz7L/DPxR77249GV
wz6zE7tacVjMOMIKlR/M24LFPK99PwOoWS2iolJ0PhZNIlhIFF2KgiEXj1SPAHzz9G6Kg3xZhWI0
wyCCn/qZxZ43dyLho1JhysXhYWRuP0hPTDBKFMX4+j/R9tSPQAJo3jJd4+aZCOPBxSpt1uJSy4AF
QND5N+fwjQWlBsGnO5wKZmMBdWYzZDIRrhvCHpMS1YA1fRuN2BnxtYkUxPY0W/2AWgl772c9F6p7
Mx22Y/91bldcCTWxGYdtmDFZ12XeQpPu2y37HhbVz8ZRQ84qzsioTSpdh5ozbyJyOo6Y91b62gEj
0HGGGjlisSzyl1jn8cKRnQYGzI6SkmDJ5XOpnGWpXNQWCX9GExXWO31XCABL7UmwsV8J3chOkh6M
VMyeDPMblgY85zwmZMovbq6fV6450k3jxRQYBl22y89M2sawnyKlH4jRWGYS9gSs7W/4Lzpldf79
kp+NFZ0eZKqhgdmhA13HXoCxlO60vnsiFvmTdX5cITqKIednl5SxiTZPBOedlAl12iaZ8/xLjifo
ZffLeyj6HSxhg4JOJ6LHCE7ciq3z1XfmVZW+dFBV0nFLZeXPoIhXrq0SIXQdAyq0upJuI9G6e/Nj
MpIuY7wREpZ17Nqfcf1rbI4dbbeaYUHwlxvyrMpo/HozyCqO9YXL6I5KURKnUYqn+oHpVt7l0LhL
C3JslyILn4eRs85TqyDBfXKPjFVQQstAmDcYXhV5ijYnDsYA5E72SXZoGqSZe5bdoqAFEiPtqDov
MhSvcHlp596iuyhRDlPbLBf1Xni9xTmNuml+/H76YjHGqjJd1xTcyfwqJJIAHnUUu8wygMuykO6k
C5h2Vx/Vtf4eyKjJ8f7zm/jkQJgv0a/3y7WLy9KlbcZEHg1bDf8haW9W/BZEIM2fzmN9038R/SED
9N6/g6pYMUPFhkeGfZHOizRNbpf0Hc1fU2YnN1sBs3BvKHcpoQC3AuPFcppimk/JgH2NwqebNf1x
z4R+WlQGP7OZ+BBrMWfzAvX9dhFDS/4N6ZGBXC3cfePkgmZErqmhKpWo3HocmsS9uTNdeBqykz7U
b7oQki+cTiwarMdEQOt5CLORaoHbIexgLcyI6oNSVs546qNj76vcLrUVby8dWA4yS6Ox1Ub/OMlM
C6E2uMmYywYWMjrFkAUnZ2hRR4M4eT6pvZfqmaNfzhEZ7orlhbSZy1XfIQuD3N80uUSV2YB+5o3J
1sBcPv5SL7iQNdCBcycdulUMyScf03VvrPxENIWvuNz4z2tFDNLpc6PK5es6vy0qJgVYNw5cJTgz
eVKGaKeIc5QnC6tCoEy3fwJcmJWtlVUD6VQOUSDutvvGQU+J6kNaeBCRWQYWoL81+00MDL2Bnhrf
R2rsgENhZPZYUFvLbrBGP5WePdFvbNpZT+5cwfP8yTJJgnVIhG/XRael6NlwmglIT92aU23MY7Bj
6M7kOXG+bYqD4rfv98Kt40asFnTfGZ0hmJzemEfd+JNc6KCWYKAGJ+mt65nvXwR9SFn5FLL/JEy0
j+z/57nl23Z2dYvpP/hcsUuJUYBjZu1orNt03uMFspajrF8uH531NbfOwzbpMtNB3X17lsH40Otq
Mtc8PiLJ3HYZyRyF5XmiWH/TsSyfKOVXMuvB0WgowEMFudwDcVAkX1OogCAIJXwex/BqdjaZyQKN
GVBgWnwEepJN2Y8yn4yoLpYbGoJExdlnzI9YngJbY2CWJV7aCTfweBQHioBDdhsETVyn26RY2yYt
C1Qbw3GgtTHbZ51VA2Z8m9+FRG1Ud/bl3usJtd3juDHtxdkXuGeGLj7gYUkHiYvw+yibmBjr2poe
uJ9o/lshrJsq+BiOpDseomBmLa80YHS5IDxj5iUVnHmI00bBWodnxF4ic8jvasKyt5y3GUmeOrDj
5UVhFkXLbK8wm/NWkZ2j2HzkR8epv5Hd2dByMd/MnBrQflnYiqytd0bCkCl60YI8S8gV5DnJvkoX
XYoFo93QAf8h3wss0eczy+P4qkvL03zefQWyDoOIrPKkkdv7tCiZgIlTIjoTZf25irHvkyPw55HI
+OmQIYAEOxqne6tzajlQs8QL3Ulk4VFUYOHopdqUy42VzcQLX7JX5jIV1kkSR5/BrIaLeqSv3Byf
E6epaihpIaWo32juG0XKBSsU9QGt+rwoUF428hxlJ/pc+bE2IitmPkenlvuHh3UGXdqO44w2H/Nc
M9GXMLmzLGfoM1uTnl64ojpL2/MGSO3XqZO8nKJ4WSmKWRZn2dKMKOV7LXciqsq06emQ36C4ZMX2
h5pATL+EvB8IBvfU6jUHXzzXyurUJMK+rnBCE6Av0cIZRwX4lPLxa94ulFbjBakRaa2sPYMZzlr6
mHg3l5A5RDUkbR1i1ah1UjutuuYxjC/VW/vonp/gqAun6l8SFFcnC9n6u1opMMF0FJE4W1NoDQRB
y8RklQ9FJOw03dqlzBIYk2mkbgqwxxNi0zN67QO+kYbE+Az/1SAU/1csRucMpUYFI0/9iaZSU6pI
ZmlXQ8FeDDKv6D+MZfy8S/EzhFsr3njOW+u6MJylkyNeWiC4ywIwHSZiHpbinTmgwdPPBnD27S88
x8IZL6zonrs558jc0Vw1pAtYmxvHnZ/CNFN2fQ9ZBQYGG0pgHKskp1bjcIl3IXq8+JnEUv8/NgIR
EHsLMgEXsRpGhNDEHGZqqDzozf3fJpVFKiLQF/SUB8sbjQyvwNCHQKKZVvMNWBGz/mLsft9B5uBy
mOPeegIxoEe/v+kiIFcnktFGjSkKwUYyiuMLOrU7YaBuDUW0h90pWTL2Iwpa4WIQQQSbUr+Nubze
GjUurVSnqY6w6b1dZuIHwTgv4YxncwJ8o9CcBhINCpnwRXINy5X2BfX3KoDBhpj91riYkXaV7Bfd
AffCsYWPUcQP6vpmWpkepaj2pPLpa2B2eWFDdFQPXQLuSiYBxXUWF1XoU7poIZn4n0lQTfHFmGHP
T0kiOy38GViT5qPujO61YRjN2/CB8KTXhsg1z/xxsijLtjZYtsZ7QQnt+svxDgTlOU3c9j6ER8K1
IwpjHJvEqKO7vvjivYQA8K0FAPrnM87/b+p/hRccDmzO/InIA41QyYZ3keGfuy+DAw5EuHbNo/6k
DtkMgNi5toYZ8fYx8dFy8tD7UYscBXUjm1IgpwM6rNT4najhGKUSQpb1cZGAv1S6IbQogZkXOKII
llxcIIZV7qSeTUGhLrAI0cdWzpmpt2r1KH5is7hdPk8aSXM94UgA9Je5bELSOg/Wahydy69qUe0h
0lVGXq5c6u5qVHG+ZqFgAwOM6pkGtL35Tb0koxnJE1fbHktKen1qM9F5BAPaNj67G9bqG7eCyMgw
ccETzXFff9+8Kp77i5f2FA4q6IwFFk+qTkPoR1eVL8l8fBAyCICsnGclI33IYq3m9VKAuIgPvjQw
WKt3WsNyVRLeYyGZIq5JiPgNVO958/NFGgL3mT59/3cQ/NcJqS7fKy3mV0zmPqO2Ln40cGBD6uv2
d5hdSRjpRswhQ7b06GVhMc2NQ9gr6m+qyQ+Nn/OEk87hPpPiODkskCq/d7VWuQQChgLCt5qi79hu
BmJHcfEH6HZ4KsPaIWTCgDxHVC62iJmnmuQcZsdvyjLemi/zqoIPQzgzRQlBkCgdWI5Lijbitfue
U+123ejzEyq/oLLAvptO1lFHJP57WV756TIBD+nJ26qtpLZPIMjIpGSmTPqLPiXOxUFRKFYwEpvD
rejL38fgAhxiueofFuc9XHi8ae1R6mkR+SOdhkHXsN3eKdN+kb2MwynSLpyChEttbYFJrdKWO+o/
llQd4zLpUvm2EysWDGysF5EkZvCejm0ttlb+C98GlS0A6YeUDAgNFrx/Tj19v6MrTGmKqamBX551
9zkrYiXaNmvY8Gv0dr28L80YLFqrhmmaosEGZmxB3p9B7xYdnWd7Js0RqmK6qBX7LnvmjboDSZWd
wJcPuAayOJhz2cVF73YfzJ3nKQ540UrNwWvLa3c8BgKPK84b49BxDwbzd5EAhwRt9PU1la430aH0
/INARz2y/0C8k74Nm+jIjiXUnUs2Ze3DpFzjDKzO0bC5dWhgp5mJW5QnlBTP2Nip+OOG6Q9YCvP1
C+SzwTtoVnC5dHfkX9YryNf45W3UrX2q7PeHvzZ9TgzHPUMcjPL/OOfNECjjTS/rwYAYXWQ9Ve47
L3gsYaP5wFd/kzaliqzjSEInR0V91M9xAg7+idIEKQPdWtYQnIxHWh6nhs3xjKZyv6mUk6NLIzZn
sLvPSB34AzSolBdaZ+f8EhBnGhAVuYw+xov2D1uJ1VK8irlhupph0WyQLj+ilrWIeRiOgwFOif5W
Wh2VIQ07+IeSN8TB2fWqYhW0V6f3quurB8H0Xsbs5rsW/oUhwgGJN/LphE76AZJpfjBVWm1M599T
y6oO2jSWzdednzu886G8TjrrZx2xdwmz72EC6E1qs0P/J4bFnRn4EYBdxZRKy1Th4fjwlF1tcM04
H0DB6HRztz9C7eHKptVY4X0tbU0QrRUUTmVsy5qDzTtImVGBuFCQeeqySM3+KZJqo1C9KyqJVTPf
Nl7lsZjMlTvq6o/GmV678SZOeXESKQdlvFV7OSpRrTR7qlHqZ+bQiuj3l6R9kKA81GruCstKGfW3
JmgAbUdvWGAFDCiWID06YOFXMPY9lg4EnlQmPZgOn1aOM1mARllxm8uVTMOfMYDxEo+sAH8H2Hsv
gDbC+HxgWfRU9XxAigXs2L8y3ESuggYR1jPhotpdDk7u53oNoFlwKJNOXFRs+MtuYNsBPei2zF/r
8g7Inzi2IKd005eeZxrdsLyKIi2IxcLaLBWRBQdJom+gSYZuPNwWIAz2oZ+SGBhvfBCfwpb7JeH7
E4Vz6U/r5mn9/g7BBVqr/P0kMRcf0mJSD0IBPKuQeAJszDTXsjaFoMj/zgRjMGJNx9yxBw2yBy9R
/Lprm8esosZlRhkLfBY7zUzX8Bxifie020y/GCGBbuVTenqLJwJpOQYo5pAI2IMCgPtNnaV//TdL
JqIkkSKQ49BFB10rm1/bUeryqcdopjn06gg3dOHoGVP26OsvN/47hLdySIG/8G6bpvW0482o6fvg
0RSoyeSYLj24umtWwscgFIK/PD2Ah1oKpzOsEFxSjyCz2WMB135jIZriKP+nvkitj97AJX2zrCgI
H/8YzokbiIUOqtaBd6tyx6DVMJwlbYamVb/LqvToYAYsCXBqBewfRTTL7h35c7zQ99qsB2PcE7eu
B+9znfwYP7+CgODoiJKzs7r/uq0vQraFuK/uok9NZwwNoJsl+30sKmHRJjOKJw035ZQ5Xj5GspIc
f2RVBOQfzawzkPTTv9Pcg6/aLw7Jr4PS/+fFs/is3auEoJHFRRKZyD37gj3ddO1fQb+m4yvYBldu
LdenumZUZFp3q6hvlWRhrUkFQ8oMt9xNG3pivUkbjlf2zkbaG8azrfj2CWk/4z+JpFy0QfnlhFHf
CfmkYDFCCcQH7i0BS10ZBI+duA8li+LBmGkqtVAcbjA47x8TJAQcmAEQMDoaD9Ch9/q20B0bixD1
R7ZrX2lJkphXnPL5ni+t3oEwBgY04l0fTOT0+RLEHa1BoI6/adpDssFVqJdrWpkiFl0t+8zm4t6r
rZVlGqzO1IEXN6wT/lIjAjFtZI90IzmGO32asZzueagTyP0X/Vr9jmh1Jaq14EwdwetJHxo4KcK2
7nJ9Re2Nuy+JR9mlA+U+RWAASS0Dvkri3n1ViZVviRaRXeYprUxD6oDEa1yuKCxaAJhQccaTwRji
XMwLdiurDQCPTbNg1k3+voG+zhEsXVl4whp93+T4SzFJas1ZkwbZnVaZHdUe/q5mCzDl87VefAGK
3U4FixyzLkwoVjLsYX+6uG9toFmwK4YVrn+j7BZLJeqBN11i8HJUAnk8t+mn45t2SC8A//HmSs8X
FBK33bel211K/e+sar+YGucIFDZB/83jMrGN2ktxys8GjiMwuNCYW37VQsZAKMtb2jrqoh852qlu
JfNm21+MruMt/N4DgB4sRd3w+JiIihCjlQp4M4rQRdS9BQ08opG1s0vbj8R9+pS45CKLh3qZd+1c
DbXt0IP4k5fxxcMDd32RecuXvmZ+33ofX+N5esEhNwgsA8YSgDKdNm7TPwG4sQJ2DDpp54iuDg3b
kBc0CwRWGhL08HtrzauqrIpKzzOy0/qNvhYwBYKoxvuCPLV64aA2HgeZwseWJ4/VvFBJGZQK8K48
j6r80vICl7zkjDRcqyO88YIPwVP+PHKrHS/FPzXLM3t5RBrrBHXL7vJbw7mR6b1GBYYE2o73Wgzc
/pPa5e3TjiHQ37M9AjUxGexVsh1ZO3v5hfvVO2YC2yEgMoHJ4ayXcuc3LE5reacQszg7Y5y1kNga
pn2XMHlS8pHVOZQQe/lt8yBTGp1O0cf+cbIPBf2FFFqfKw+kpV29wMYJjhSO1ZNtwV16WBUYh2b0
w9cP12n42q5TsOsKmmpB2x2paMAxnVtrJ9wEFcWHTuNneHr9bdh8i0hV0t1lQ+TJusleaWPSok1J
u67Jjax7dQ9x2hHFN1ep/y6NnObYc5nmFAzkfORNw8rkM1d+9BlWAppWPMoSvKcVZjlv1tY/QwVW
aF880b3k3s7FXUisIF+grheqmho1cJl3bRoNS7FSsuUYGbnTi7GZtRGH9jR55vXOTvIwF8Jrrmfo
xHs+VqqJ4jnaMgn2cnBZJx9QFObd1lSo+yngTxIXDOwByi8vN1nrrZvOHoxswx43EsyhXdWyKqoO
D20m99OKuF5vp//LdB0C5Mq9A/v/VodrknaYSSGbu+7xepJUq56Mj8jifpF2orJosr9QP/ofe5ts
3oYGhi+cLEVqas/iy7LW9v1JfFinGKs9Fkc1Vf4uN155/gPkNjEbkr60mfsnDxuDovsGTqG08Um5
CH9mj1Wqosq4gn+M0eR4vqRTTBcx+o6rPOMZaLSl6wgcgt1GacxtfoKzVcPuMm4QtrZzBV/LucGZ
SO6T2DvrwgRNcVCiC+/MZ+Be3Ef/vK4aiIfZ/jrXhcdleMM3VAsgLjIOy/E3ySamyZlPQBhm6SxV
pnkI5THkTYDM3vkmwKy4LA8RBVSEwkgQNAcMJOSolCtUMJvB+5wP+8VdBLZkmmMFpF/2z7R4PjAP
jl8L4Pr3MeuKzMPHBvhJix+zIpQafrgUHX2yZf1HnvdmzoZX4nPNLrhAPtjkxWVtbUWFYbYz2DZO
9acnHaxEGJ1BiR81y5Z4AhxePy9aylI0CDgFkLCNhUc//Y9Z42uBHWv94COojQ/hgG0ZVgkbVydi
/bgwe3FvrbZ0hNqLx8GxRIFPXfW5sTzLjbj7FbDQ4YELzI62MRaU9RkmrfxkIk+RD1OBtAQ2rHYi
cYUBaA8PySjgGODDcGMZ5/gOIeV4ZNpoyngHP5l7kshwV9v7xkdTH+nBfquI6iLRhAnNilA25aN6
qKaAJGfrp2bm27/0vhjfN/JtjmtusC7PNxWIfdS3FnTCT2azAXFIFpfVkHnYg7i4kNHnac77tjk9
jNCBuHD+GrZg0OC/6BGY7kFslIha8EWqk5gaTpQBTCkEd6Wfngi4dUa9tba7AOXwwJlGnvx1nYwk
/c8UT3pfxb9op2XwJiX6vQy6crBFjbHv4seqc+1/B1KBenYEHHl509iOMIKyW4eONw0FgsZxYsYD
0dmblmhtgAkzK5aQTeutxJbSPmlaSzigR8rDBar4aTGpeNjZtQ4vEcchXpxPavqfAIhVsABZT6tI
mSpWMJ0fSIwwPPor/BZe7SGo7Of0fC6CcNOD5xoV3UnbiMNH0FB3RCk7WBuSyQKJInnzouyMs8S/
zwGDov6/1ykkqZ9qNF6H7m+N4kS7krrfyRbIna1K0fzGe6J6OaaCKRnqJsDBi5iVyj4s3bY87adb
sfDGaylVi8WNI93H2BLsVhrNNKLlUHJGdzF5UIXa5C/Wb/fP+TJcc1kCFomqg9ZZDtezpBxGPu5u
7YqvbRQ065EU8sqjCRc1rTNjvR5GrACbASflwshcao4VJuXUuMYZwcqtFvP8ugelb3E013Yf0EsQ
ErvrNvDFLyuLafsrAUsyqeYQC9PJmc+08LOlovP4BGAVVEHGH5PxgkkKRXlw5SczmsWZ06sghn0N
fhAoafoLnrOywdiCFP47EeX4RiwwXHlyfAkEs2ixIY/YbBHD6I+Nap9hAB8ExNQr+3dqou44S94l
QYP+mhIuOi75rtpz+lHZW+0o3FtONGl5DMdl3SndjqHRydp1mzWBF/QWG8ojLp0gRwYarLHyP7tW
KabwyfUwrhSMOZpv2HhQD6nZl3gG58yBD/gZXlVcE76VOo/EMQCo8OonvQFOAZpUfzY/NuoezOA/
l4jCv4jqmxAYtu0WHDkJKbMRwP4M8tQ/EWrTfVizwUN7DvQ+3fNvSBi+rhQuEGMJuWYh2BCWDd7B
3WRbPHUPK7d9b6E7/6tOOhDgPA5lomgXPAkBzIC3XAljYplm06GeFMjOzp5C9nbeGe/1nrWwkYLn
QJpg3blgJbKzEtHxye177Fa3Z3YNrJCujfjk+0WHx45EtOI7NR9FPyFcwaSnLada+LbrJ4gaoTlA
w6Q1YPHTascVpn4uslT6byVfoy6qD9oWpgBOGpfcf+aZ1T3USmoxa0hRfYBcv5btE6L/jSnd+Bd8
ac7x8Jg1tOBD/DACZfaGq/cvgrqKbtQ8TWNmNP1nA/iB3h/zP5+dWLtc366LURqduDscnfNQGfaM
CJfDKBSh6++tFrWB7Dc6O1cz7EM8XtknEeJ0hQZUqG/G5KdfWnAMzWrel+299L/yYszOEgSoeUsW
JZS8/Aq4ZbOb1LTMMuJLi3lyJ3AxFPPeifsbfZvg5LEfXrK2AWc0v+olkSjDqa1EiAS0vpe623lS
ZaMRfufVrYq9Mj1bfxRwbyfVKpKge7O4lidwLBIp81JYpGdvlyywMIEav6w9or8+xlXoEP4tyGR1
cKLo9gFj5XVdL3v9IrzHNMfUyjbma1vNCbr9R1PaP8JzzZd6xDJFqImw1riqDU39vujfYLE3tvG3
rBNKnPPl7HtqxKuMcbOwpLLURtGh3mkcayPZZuRo+NzPNty7N73d7y79QyhwFJWkMWPlng7W/R0W
z5KEM2WS9PWuAX6Mtm+5cTL9bxS2u4ExocKPRBTuDq8GoxccvA/AzcXvQHfOWQmgomF+6/gR477E
G4W5CWxjHWJ8EUgvfuTvPlBfUfmFMqfTMSzGZj2gPNoJRsWhZuljYUt5uy2bDhHLm82jl9SKrnM+
YKRzQBCRJc8Q8o72sFSrUBLAvjUkeVYHTRHM+DK/Qu1qYQ8ubEw2Kv9zPjLZAK8Wt6JP80/wwLc1
ZyFwVkLGlfNOZzUBv18JxoOFUg9E5OzNApQPOJ7xWfFFOYnk8Al+5cuAbfFIm0mn+CeqS7RjWvrj
qjUjj6gkQsiHvs6bKWoAMDXR58H9SG5KsLUQRKpmc2TgKS74VoZFRHy5OScosUiEixUL7ujbgHVW
uccPS8NQOOvLO4bh8cv7SsszZEsu2S8phxCreZg1o4NCiiC5StzzgZKNfIpue8ZGKoZM54Bw6gKx
RQMgx2pU9Qdp/wlAD0A63qBwcY/moe9SvlXArOomzBEqbsN1Qj+jOisntmhsBFzbHu98iSnsflF9
B8ZZgLMnqYtiewujZcf8OTvTh9QHAV6CbNlwVCqDkVEUUXC33wfS+TaTLNOObnrlP4J0PF1awNRz
AKSLWL9mlboDAsT6OHSi+40goYQQxo92jhpRYMk0xdYICFrvw5CB5ZjSRU2oe3rbXCanWsNYvYHv
lPJMhrjH6DWESLYNzbp0ALhCYR7e+8D/AIMckOWmqkWn9lCh/GZNPfmY2O6d1tQ5mdDL5JnqLx9o
9wblTTB9zpZhjTyBaR6cKn7ynfnHT51zmqQEnp0GtnQ2b9pPu4ykoXv3XVeZmidcftoWTmXJJCaF
LctFCwSqKl6Q/9JwOUzvdU1IhwsOWxJ+qZC5xuc0lbRvtZcC64XLF0cnbNdYlM/gRUfXpagxphaS
qN+MR8jQfchfK+TeWcHWVtMWtm5nkC9QVeWLrm+h2MiwKsNJu6QFJDP3EYG9BCYijV7yrcEcoh4I
xKAsgHD+94xDdHfnymv40o8oMdhTcB1b4973dH8Rt6UoZt/BjczPo9d/rW8tCwgEZPfuMCu5o4qT
7LDOZUQErxIzb4TCKHIjZ855CQPlR85FNy48c2Ph2BQAkGJ8ziKe2FuLy11gfSUcDkE+vZVDYYAU
rl6HiL+9CB8jJNj449h6Ao7yLBpUvjT7xDIC8Q9KEq2AScNh6z3jm+p/7h+WWqf2QzIrywF2rStB
CUWssqjk549OYEPpjsPAZI3c5F1P8PuZwsAn4QDE6wRhE8ZygGXVSlfl73mMkB5DesuBBK72nlly
JKb9IDt6d0ESt6DWoHXzO5dc/fwQKQqf7+T5Tf4UtIqK+b0lpngIonqv1Z2p64Ojt/qiqSWii2pe
xgpi/WtBdZaTxnZuF36VXf5NTd9KFxW64S6KyT3aRarQBCAXfaVyj1KYoAiHD463iSWtIEivt0OL
y0v8iASndfo3r11D7gNdYxwE71cDMJVh6GWKj61aTedTaf6VUBk007btJH4vVfejh3DB9u9qY7oE
tqQOcfyIposc/NoZFkVsWK9IwV242NB2QDrl1yDmDjUK9qz1dy1oUoGZG1TieDUn/RBKIpTCpF/d
vEIFUq9d1SGN+ohJqMOxvtx21NrXbu/IJmgEfQq+Wu312MdMnoSPBGNvTHK0IikVC+S27fJ0JVZy
xHmpqRKjsyKoEpOKByg/yvTEPqFa7y1B06ayI6gG+QB+a79O35k3UzZatH32L4X4/iIoMiCZDxGh
R6UVkWPNhzsRHQ7ADFXC04ZUTB038tlB9MD/KqSZ8B1bRemggkeREoxo/ZiTGX5DrFsDxjblScnt
mL72HlS+IQa2f0NSoV2pvyAH95RrwDfHlSn04JeB4AubUDUCrAEliOID1nsdcxLRCDIkdlSLD7fX
+/rbTHEGTZNTvrVUU4IKsVvw41F3ht/cHU9ATUCXoDsthPVsmh5+W3y+6F7O3em1n1Z8Jg+YNcYE
wuxdu0xkixPz5ZhNIKpP2YgqyBqkJA3Vqe8a7LBodKV+QUNaOtK1/7wcnLBpK/CYwItLSzEfE2jz
1dzmTtGei2Gne+oIeS+UyyVAYTXO5jsvQTDW4W4Wsoyz57GxTVyiN/2NBJUpZG9Q9t0fnBXrWX4l
cEJpS0BwTyxCumBu++8cMtratwrelkjEzNu6kdcxCyy4gSxm8mo3S7rl2j4g/nqd4fD/kvLjQaaO
GYoHl0y6EyNdhb/bur2S5gBFYqN+HN4tTpy7otIzgfQQsCFm1lvq0kRXaG38670Km0mF17LHkogY
qYDFFgShuGh0hzq0alINcFrzu/OTe5inYAhIfyT+wqf/gcJLRkGJQO2ynkbSb4AMX5mwtRaZvlTa
HqmGbJStUKzd7Pgbnql7E7BCUAi5bX2J/IuojE0xMgFWEXrAKbmDxDfyMk7yOXj8pdZmG3WELTbL
RTUsXF4kFZ2z0Pmh38EejT4A85rSYpWBLr5+6ScJLaGkCPSgVzUmrkg65x2GDhwL8ezYij78tlXk
Z11p8Or/lckUUJBtEiN1vHlCQM34o+76v6dq5CxUdKMiw7dpwsQehdKftxWp5ZcKBJNlEz4aSKTD
tesX7Bgu6q00SDN3xAWZ77HI0ajK8/Y0Uzu0cPDfTZANDEJcPVha+48NGblJroWo6uxxMnkr1mv/
fX8MwbbUjpR6Ab8UlZkBw6gTWRJ4Ayyc8GfqJkQN5j5aAPXV3H3Q7jRraMOglA7GmYexOvRYjgrU
5UFEYc9MYALs2KmO1MCnrUoAKmQujOCPAC0wEyuJjAu0BKYjEN/3qyNHbNjBoTk0IUqUy4NsORAp
6bqFR6YOpkt8addWGYx9Zlg/biCGQp4U14Cf8uO4sVJfRvoBzOOIDPVWu6eGpskkr0Y8ZK1p1v/M
yElwJ0FwcqJlhHva/dtK8eCx48YOSQcmYIwVINuF0IlkABVacbs2S6iCmL1qMP6wjTtVGVwy5LGk
na1hXVtg9raDGIcihuq1s31ctgKIgzXJksvfnycxMchV7BmIGJcvEu2TnpLoH3kNgvQFAftdlrrn
Kmnm6NAQPFhYTlyP6ZBqGFdoXn3HrE8hTrAJutd2SGSb12WZmHZhDC48Sw7QFKM5Fa12hzld6+6G
p/sPwGSp2nUG57NDmPiBMYV47gOblpG1MzKXHXJ/JCL2ckXw5PjUlCANpxNMjf6R+taNNSuKeWOq
8UqGnCxdcUUmAX91axqHrRGJ32g6ISjUUQxNz21Fw6j2K1nHw7BRfMEw/l7fHIHnpO998l+YCnyL
zUXBoPF7kxuRYanYkf91ABE5M1Pns4r3H0Wa+S4P0bb07UsdkKTFLP8FO7InS3el40GFtRI0o3DE
hl8rhafTzeXN27sXN91n6bgAoMTpwGVQRl+lwFImHfg1s7OL8d9chhK3OC7cTBcRZSk4BIZxYpoS
QX4GPxPkW5fxzs34SxKZdm8XHq419xJH7jZK0jWFWWwPCq/WTfKrDvY6ME2C3A55EPTDr49WmNqz
hXZFpG2NEEZW/HO2t3+oewjKUnFv79QbzC7dvUiktXD3NdDatBUKaByp4irjPVn/Z5KdOJFf2hue
66tRCLnBFSIeq2gpkHNz2781f1u5gTi1ov4veuuxfsa8uHdWCuGkR2a/SyAERZaqPDD14dlAGkU2
I8iBaJ2GgOSO0cluI+Q3iM4AkdeNhniBiad/t8DDOsSzmo+XOC1Xi7B4Z4rScp+DVz5g2H4Z4I56
VA5eWiPZxoBsFjV/BsoP/7tJxtfLJKejpNFWuf73mRH+fEBD5EwZvpsfx+AiGDZqBvFvJeEeOQPS
AzzVE2nUxbc7cp6z0/9M6Zi6fu9fvU+CsSshZbBEhXeks1G62p72HOHKmCrEARj9xqJkIxTnpdu+
aLwzLWmcBeOcMeabB4D1B1QgV0kJ6K+GJM4iFob41kVYQ9XRZS6cH1YsZVV1DWw2gOp390+14Z6z
t1gFvlk7EteZYQ6hJLD9FD3cAqbMgWmxIX+1B+vuSV31wRgXfaGFGei2OU4b/LxmMimwKQCoMAgA
RhewViEQ4/ISxaXmpluNavKTHB2I53w5w/lg7OiB5hvqv3up2vZz6HmqRZXsW/sgf+ZkUi/ampha
f/YEud/o+75StORe6VIx8zkxZyOYvxhKVrBOmpMyegUzPdbXA5ROhNjXnoueMi+aOfqgZ581TVMu
JGXHZNxMxTdwXgHz2rXSQqny9mtkFn9bxSehCl2seM1SMSXch5ncc46slO1MG6FFhzzeOUxW1SGc
aD4k4FR1974oeZpkP1dQ0tbQqKPeZ8WKWGCJJhsZaLDRuK82QAR6ywFd6hYumZH3N2WRk5Ah7Is5
aON6108qYJG57PjaGdqH9PDKU4ADR4jEycT1XeOYCmKwmUSJ9nJgmRMqm29kS4ilAEot8+WBz+Do
1evIZ3eDqzcK6j2xLJ0A2rL3to3eW6VrZf5URfMDZ3qFbxXbyN4P2vpbpDor564euR4FNrTQd6sa
1fndqb1X9KZuIByUSz7hH28AmmQ7N8n05nuzyXWZGfzrXUeJRRs1aKmML0rATktdQ4QxTRxUR8+S
kGHeZaV20HjOr6aQiqrXo7KI80P1wiGZcqdGGZtTy9NaoEj9BAHCjTk9AWTdFEmVaqD4tLPZogzk
rilX7VYJR0ZRlpYsuQWU8fTTR8p8zyFThpMHb/4W0qA3VWHiJP4Smz81a8vMRavkZOL3FlT43Y98
CsfbE2DcgdDqjD1jKKd6MER3XhMEwR5hpNagqLOC7Y8MmPj79NM8XhiPGeEUaAmljBMwWkCDbLWi
X9aviOIosz3mFZM/pvAPYo6JfJBVQhB1G7BtLL4/xVi0JJiK9yrjNnAEI2WloMJCRdM44BoEADKQ
f3+jXfxrXS6e393FfcrhEPdbOoNr2XblgbYomzU1rjG0J2k2ZRNh8WX3JQNbEu63Pb5C6mNsuWu7
VtZC7r5E/dZX93hSpFBzK6txMYPpD4vyyGB267Al5X6qvgWRWrBNY17wfjzM9SSNjqMFQyk3ypLZ
K+7Cym4JGaTxOt2gBe70eyAC35Q+3Pxo1rdQCcmCO2NKFb+S4e994M+Ccg8WArupNNjINHfPwaKI
83voYx9uaVkjzhQbzpZy8VxBxgrYjgdiRmggUVqchW0+J4egp+1JNRobVwQYHCr4OFG02E1VVLcQ
A1/MeUH+BdUPWulDS0R0cN+3wqyqTkeozAnOmVzwK32MOBqgc/zo1dKXP+lvSEJKWU5zq2em7bwK
hr28o+tu4Ml9Fsk8qHNFAzw/TgyV2qSq/UITMpwrfXyOSIf8eDuptjGgCxiTGl4JZkPlkB28lDC8
2XUmBE5dr1EqNyrbtg1U6EpOBYp3MkD18WfcMJO8rjuFsELd3Dibs/HAFODU/RRFEIQT0no9sg7c
FxLanFX5/Mj0VkM+PKCPhrc7rkZFN/Jci8AS5SDKzQ7TLM3hWyXCKFhphGQgEyUHN+VBJxbjJnFc
yWNjZmCBsfA8ZUi6c+HxQLGEgIT92nqSKqOvEzU/qwYQHJfd9+mXI/8LXVseMhgLs2VuJ5bonm4p
OLogt4SsAT5jkcNqUVdj8JU0xFYAlYkvFx5ZBTZdXg54HvbNWq/xvkUUkdrKGFz4tmCUK5TOV0Do
tsQCgcMIhdDdELQOyJhHWfoiZtJZAQolZNASJma9ihVBQy6MYjrMaJKzwvlznNbErctDiuz9DM0r
NGAgjFOXvs1TRdFil7NiazlSGkJOKA94mxbFzSM45tnHgFj9MjzojOp/fBd+sqg102daZU3dOW0k
fwFi7U3UWDN5OitbyEHyPe2uvp0RcwxI5ypMpbUrJQceplki6/QccCXIm5OSo7xdhcSY0Eq/fCne
K7lzZ4T6mKlugSkWvYX4PfgJo6fDfDzGMZMMnvEgEJhnCm7Zi546C2zz7oikJrTyUAzLbk4Jz6VL
syyAnxZE/uZZvHcHavXZbWjtst8vRtuXrpTLsmtD92P2WdFTcNU8GoYpLiq7q37wTU8tqTY5C8c5
poosiLSECz+XgN9t0lhaTij9fl2/usq5pAG7AkuB60bKpPlOVK/AT8WMMiZGhvuOZ4khAvd3fvkv
WiIstKwjKbe56zAMWWA1r359QXy2LUK6EzvTrqv6oY4pTUUv/neNmfF3GBi9BaOzhODABi8axr9J
3abz2BiDGIPze57Og/jjiVYddAOfZjrsy6hBN5ruWVqOrEJgUyAlsPoOEo/YlTkIJWT/F6yGOO46
pZ77zN/Wl79+hR6qBxpE/r+cRRl+cVanGy6Hu3cWAdBZA5W9IX71Is4gbONCSBrpl8lLuldC1g5i
anTCznivzF4S5mgQq1oFFXFQq5FrBF5y6FLbcWokyexPuizPDdfME/Bj0uKfG6LbN/n0NOxOpp3L
hiYzspilDDOYgeZBN36Z/TLLF/HrputmbSjLv5lLTn+IkP2lddGa/vx5UN+QW4ZLnQuRKs5nsI9B
qKO5PElwOrsSXGjxFhY4l0ia1MD7HbuWXPIFmaQxJ+MCUe2EoWxdCFSsZYoitR14EkNaApxT5YPO
nOsF0Uwonvy98Fw5eE6p3knaKDVN4p496zUCAC4JK/UaM12oPPZ4qmZfiI4Zk3M1i6H1NvQu5BkK
y7VRB5PWOU3hgyiv7ZilRDKOe+k1Pg9xoRYQlH2pBu1hz3dCEeM4/77jEW23Z+0mI93pohS0XN2j
Nk9ZKkhj0KNYN84w2WBxMpWyKuG3yPoDTEdiXoGTsNei63hVtccCSEGnn3lcgtpJ8VVbe3PFAbEj
YeVc8WYibfCw76kh2deaOTD2qlsNnqCObQGlBDuqqvvLCPQCoOwCNG13hZC4NCkihBVl67j1U9tt
K75cDuX7LFa0wxW2k3rEwE1cU3W5v+htr2Kk/cTrZdfeu+ogmDwPmpTQGb9PcLmtra6FoRG/st2z
/hqTMPk2ZsgMV8NY+HiJRTp1jhePeDonrY4qP5o49CQIUoeALW6Wj39lQpAe5GaREbaInqyKHBlJ
WeZ5yXuIukDssC86CtYT3ui1KvSfETD0D5MzG2GWHH2pcAmr+ie9tlYrKAujTgeUdvApcMsATsxG
gNQDpySHqfOQ7d3knGnT6zejeZ6gcMfees7AP/pimbdFl2bo/s6xxv3//OBl4I0RaKo2y9YvbtSB
LSe5qTdNGrzoxAS/0qqZjn8CgHGgUK2ZeOhxMJOmxDb23iMwYuxHmOt/HAm12H8txpNV53KvFP6l
1AlHxy8qFvzme1G9Ag+O3ur+F3i672CKI7bNrQ+Q2dQO310Y2868vzrW+IMYKnE4JwBomgaTkjGl
Dz4BI2iGRdXwEO/LdcPUkBcXfMXK+UY9V0neleLdYBoojQz9KBD0mURDFRhZvlKdQGtHJsFVRQWe
Ew2DvrFYymhoho8IDRHNve6tTP11i0OkAOceNpeKDLPtDt99TbHGUzgWGSP3hFdu91sbjAljYhtw
fadYsCprb70vXwHuZnk3XljOpK48qelaS1sriB8alIlVlkis7EnYTGOKNDRmNjVmpdYQCVslRz6G
NVahg8+0a8XLzy/musEngdcEf/tw3hJPh5ZDOVDVt/2S9dyIrTdrcZ0bPok5Gx0Zg0fxEcPRrh9b
FOWpeHHXd4hFn8O8ZlarntwMQ2K1YDrxRBU/qIwlsSLqtcxhRbUX1GF/HLOFHKz+LfjGTacimBsA
NEeZ12VSPw+uo64FQA0Hb4LNDY4jp8AphqTkK8JefpyTeR5QIS+FzDRXhL5EdBw5NxDYyQQJDw+e
mTVxaS9VOk7TlQPGz2A8L5044iWRdHcwMBVuogo8ncOx3jFDKFCIvf6/EVRj09SOtSRxYJAlZmcX
6NDdAzCpLz9QzScqvOiLqO1a01Vq/3BhHwXu+ngxneKt2WRUJFDzD7jhxDfIabIIQ2Ykdl+ChKhH
xDYUse4JFEGyCuLbKNQcoSOyiahkUSNuEf2orF6J11aDOAH8J6Rtwv+ZVGPQWz2zgAZT/tPbNKw7
loaKxjVnagMaIqrdO/duNjnCLZRyRrtDQAK0hS1oFwrZU4U7IrVcv+MnYO6eTjW8NWfMZEBeZAqT
JsYBQkV1rIq8ZfSR8tfRFcr8XNggeawYSSLo/5tW8irAKxUIQi+bh6NZZiJ/iHiteh9/V8Arj2up
djBw2OROvs9q6+R15psu7CqpFg9yP1JK5i2RWdI+g265hmRCzqdapJmF6m7uyVH228t784lxecrF
sHrM02dwKLl5Qf9o+DzcBL48BzbYLiC8kuTxlGe8hZYkEh8Nttli4TDAbeAB7bGdrhNOMDf42hAZ
wottOhz8W2bP4IVTdyHpKFmKFTvfroVuzho8O5u1t8oiNYbVLepM9jxdd0eRWSqKo4l/DcuofD6u
ycNxLoWhcvb2gguXqfgr/n0lG0MQG/SYmsINSvsCIV3EVgVHWAz8KqwKIdQOgTlCqC/O2PMqd6/a
HCLwXcBiWK/ltqYPE8n2bQ7UUQzReT2k+9Io7o5s+rAa7Mn6hGC89K/+0wWkaM/iASicgAMuBjTF
sGIJt/3W/XIBNtcuAFtTQxi6qFBPXaKUpm+3LthAVm4Jnc85HJZ9JNIKM/mihou6ZELRlRJS7zFt
LKx+68gZConNckFKTR4PoiDqI2Z0RyiyLgJrPOgQotydS7zeCZn18OrvGQMzTZEYW6lt9q6JoCEO
OmT8+XIsp5YZwcUiemVrf5YpS4QA3YMiRVSwYT1MqnT0JrTfN+TKIjrx4LqT1S5SNspbK9hlow11
EN2f04s2QauTXhdI7pKCpPeq7yPkjLwceqY5i7WIvBmqbm+7BZlNzUFpkDk5XxGyzbAvv0b8f/gu
JxPi3Vp4Oj9PiP0f96eMI1eK0P85c5d2s80yXtsF2CE4H/4Ux2ekz7E8U1Ec10GULwRhtaBGcHrM
lYemG6mNffsx2GsLQIV6XUGqF53mTPiuORswg85shSb5JDd5Jl6cy1fi14f0YbzpV2R9jGrOx2Wf
T73v9NF0gXx8UYcAl+fJZ3s22h+eBZ9ZOKBQOpVQfoUa2oeOZjhrcys8k/w6BnoGgci8QwiU1d13
8HPFvHOS0BqYLohW7+mBvy18qEl/hSQplN0ncn/pyclQfNFABZD62hXUcHxHWlzM1jlbugtEfBjf
hZ3+Icb3ri0KkI3/hI+DnKkORJQ8YizfmKT3e+380MjQD/i2ehKGJLxq/Dyab8GI/MEDYpj5WV9T
5bbsJJtlIrGlmOvA8QV4kKWOuaRwwA6VWaqpqYlcY/bRueZApRwMMACAhZ0MnfsYa3hWqmof7Dd6
91Y4UyHpc84I+fOtO/D8XdjCM4NW+NmT11iIA3kHZ/0XfK72l22h2D294YDF5cFulDp2Mq5AgWHi
ilPbYUZtNRqnvBnSukiEgp1q/EH/Nx/7wRGySEdDZAHA5IEHyGvaxW0l5BBhgZiZxUDNkrdAIhT3
YHcaKl6IqF41feUqLWcmufOAFl5gOB9IL9l7nrsVM4pQJk7VLB2o4p+yZEM1buBEca0Pl4sjaon3
Ini5dY7NhZ33N81KCXxIztJ6YZqM27JL85460Vat1/FO2dktCtU7DBFlp9HA+X0hyQkk6HtUO6lc
4kl8T/ZGhqSHmZDWrY9r1RkpVm4yy2XHDRtcjr5Nuewux9o3EJD7OePGPtyvidxfFJUuwmopuEpy
o15IIHJQrMtiRojAbxEjux0tmIBs6BL+7VlVG7nZJcr4ac6igdCoXs/2uwfPohtZVlbMKQaERZRW
bWONSIolhHtP+O9x0KZDPxk3NK+5O2M8do4vweiZeZOv532BHSZeFZAJB3FpXNDU0UCUglfRhBmi
9YJVeJiFrJDE4ie4Ul88ALhgn7atAXetYrf441tFUYcTcxo/kVki+8QzLSwV1MUqULDjcPBrVDvT
Q79c8BxDsZccY3k+coKUoRrMNebt2l4FdfxbCuNGMoBYx4dXY4IMW5t/TZJrQtkpDA1GwL75+H1I
BmBBWA6z0aUHjtupiw3Vbo3se546dQiAvyfZgiy9VMH8PFVG+pUYRDAJWrEJfEbxnK48OKx9Dg/X
B2RODWk6WtXDThxEIKqXgTFAMOT6syVu/qHxdIap8u8JQeW/amOBA+nhRq39noD1VLQoEgsRhwXa
cyno+jatDslPUcFX1UzqFxp4UjvcPrIvzuriW8hcHgTPe/Pzrpy9c9jY4BHjhkbre9Zgae1NtIpW
wQEEyeyPap1DqYEmacX8/UFoxwRoLAlP8nV24zKXn706jGQLH51LsPzrqVmVQMMeuTExnPuom6rS
H4xFDwe2ChPVfmg3SjovqWYeKsCwIe94szERrZqDI3qUxGdPwiPfUdu9RIQZxXLN4WY4YfpulwPJ
EPOruLjPCVEXLlRNVzhpy+5t/zB5k+HR70n2wKeM2QJoYLcY9EylrWQjDSboDN89IJQovhupF0mk
g3+snil3KuTYSLRZICwpNp102s1dk9GipTpVkHZOVUaai+SMhBZaoz6h7ebE2dVOwh9DXHEq594X
v8BiilmhzpyR3/ENEhR7WCAtPspsvCc98xkX+sfdBiHpxQiRmv001jLLbkTTj/ZzM/UbcdFoowNw
PstafaXcRhKRHuuqvUNLsOcnXkodS8J5cbUs6jOB4Zs4Wyr5B62GCqgYnVLnBhccQf2A1uHWjd5n
TDP1bhv+MlFgORRzGjhDw31NSX9HasX+EMF0g/L8mX5wHhYZ0izS4mmt8JQPCUCIkYLOhrPcsWbd
HumLvur3j1d0SY9UTMv7nwqYS8mmsVGpKJAhQGW2SXCU344Ud+aMxVnf31iur48WZI+CeGM5hxKT
PPggQYrlbtVYGMrJxfs6YHlI/VKZGQ4H8RUygQgDYuUh2pbtlED5aLOLHgsYW4hC/GlZy0WUf9b8
n6XnkEOeBUOlrt6KOsX4FRPMW0BjvAU/8dTbKvi4OmDSx/dGc65ymNF7nd3lEZHOEciVtqKEaBMX
90fkGIdvYsnXtYAxtigoL6KSyUhaFzFdi3P01y0memCYg+XoUDOOuNIULzY05cKZePoQ0nTMeWYR
2SccMI+1wy0D2mhMz31QuVkqOJ+bQVQZ4J+o6AGSlrImfWRqXm6PWYGx/ouUNHSFwhiTS/SobplU
VD60UPkxh67R+yQnDHacxa8UXJHiN9vdNb06i4Bzj7+kwmeSRUpfMU0PECgmNLJK8nX2cUCTt5fU
KBTvYarce4UkbGC+yl2B7fzijPaUH2gg9j+Wl5p09KIXjcf6CFNPWMiqUprspCZLn6Uqz3DjyW2v
oUpT3U6hU+4Gg5Rku9G5EPuog3RLcxASv5i8rgt8XltPBK7Xq/M2S/TeOAE9aVlUVrM+5IbJ5UuY
+vMA5e6kPzcRBlWSklJOCna/MU25TTPpR3GB2N7s8qoQPOSgOXN1afhSvpHSC11ao8Q6h4bvmYly
ojxekdd5uUYaOpStUhxcKkrz9I9Slhh+fEXU1C9+YL3ubdCJDBuHk1U6MGaQIG9ffI4WJ9atlnFv
HekyF/8gy6sBCR9gdJUP9TCE16QdyjdeqeEh9/WqZbSWW53B0K2GFV9Kti7/SAeVlxOFBubsed7a
GrmLCJE4xkyNn0OB2/PxsNxyi5v6qtLN51G8joHDVirUoHq0WtNPINzP2J3V8NKvTkPHu7AXMCRE
XsJs2/n+DZ727zVfPvuISSHU7aIleRzuuO8MUiIYAH0FPxkHDZer7fKxevqq0xB14B0t3hSP440h
raDMK/vGHbYp2OB4JozcKt8OYXx2AdaBx4XZ6M4v2PnsqNhNiXJrWvBzAOCKJ4BQjn2MtBoxkbLc
hcHgAWnv+xsrBZ63kfJLBxIqT1OYPmIgDVOqwXG5odccHgtZNGRH2VH1KCxS0FBjVLSMqI6dtFM4
PGpiM+e8Si/6Vij2rb3L5GjtKRtJ1F7Fl3dFhbnus9EmHb1YKtmqW3mYJIca2Gy2L3XbeXc5somL
iC14MvIqv+QU+u2nbeHNhdL9usIc4hCmAr+6xrICMJVCoT2wHyCcByPpwNbSskZLVDStzfgVsE2D
sC2wSfJ/6XVmLBm58Qm3f/o53Sf/GouTBXzIib87Vv7/vGYn3k2uVZNoPZWlZubWkiERUg24iOEr
JGajGGF8GqjJ6BZOlr3EuMtXuzYg28VoBdKc0OoVtfhLf+//e1K6Rogm5CZ5d0vrg3GmyMlyaruh
HryE4gzQsCVs7S31EZBtRQHb31MF0GT2gBZo12cyynQAkK6COm0dh2CTrju5xWoArrY38FrcQyR2
IeU6K9e41ZEsg4ulZ7YbRyWcIxNi/ySv2Z5ZDL+aTIJ7BzX6mAkUZWFfFM2KLdOkhDpnJpX/Fc2C
0au/4wDzqUVJXY7YZ7jCkS9lKokkVIsADTjc9qI0gvOma66xE1uNfPNowzAVvBoNLnoogatmGM0Z
vkDfcXTVaYP4t/zkMWLv4Omb7YSSTrbCNuHb64LMjD5v07OXWKr2bEw5DoyM1V2Y+AVEdD9yO+du
lqiOy5sgE29sieGzGDbFHWKE6lUnWeCy79IMOrccuWeuUc1joYp97lPQGk9cG7q6ZaCl6t0vYpd/
1cdfHvqyUvyvgk+V1ld7y7syBE8YxLReS2ysKynXNRO8L4oL845JKJtRcs/+CvMfXOlHTKqjBxcW
S0l2tX+kuMLdQwEcoV7vQjXblvtVuDythu58U/sPuekNyHSu4ucXnDZcxGqM8DhnyZrVY2YjuOrq
CZlcOgR8ydeEkK1qttN2t/y3bOrqNJQQhHxXjjnKIQHxh8f+zM+AqYRd2mLzoAn3HpACedV+RzbY
UuWdn74It4yTED6TilU2L/xH6DcK+50aOuJzWkQCfvsYSqtlSlGDfmClcq4Jd15Q4HouBypkRFJz
5uU3BT/1H9ay+HM8z3LTqRG7CsqYvw3O/Lr9EZjta0brbGMHydaPh3jZrtZAjrZF3P/2sV3LO9hm
yxGOpc8LDHIZA/vGE8bTXtN9G6gYoM3B3zXmRZ+2KiScPGCmLlPbXwlksqCI4bcVN6y/OhbhzXOY
LysX58Hsx2kD81xji8eLckurAAnqbvenuZQQM97OMfNfyvY1OfPLjRJP4fJWmcogFcdvgC0gwVfV
8kKHjwSLQTL5HDVXB8aubl9iLpBWXNB9h2vEQmsOj6AmQUdwyN/vuf/j06bsswe2ZctuEecQppKh
HfdTgDDTThysqYQXsgjxMJImAhcM9n+Ii4gnxtpUjsPJHVdvFm43LEgX1u+CUgdSwmz6AfDI4nWY
IIWsVbhnNVtoLCvdkjYMXEDtEWX1tpmM4Aeq896UF/uvItXFDekig8Oeabr4Gd8WUy5ODVschFs2
VZcjN2VzBBn6IyIRGySjqThNwOL1o5wl6kF5MhFbDvymEJZd7LjRitEjCFlaDvG74chZHCP9HMJ5
u4P47dkXkE8Q1rUYhmhCNc0mXDlkRT3hxgnrleZbG2xGwQfDtz+q3HuJ9lUhqpYiHl45bq5G7SLv
fWxYbvtkiMeFM6JW6S+MvZQKRFNftPDV4YTIT//zFMiV/sO/IoRSrrs3qCd4J5Mlq3tzcBwDvX5j
5ac7Yk5pRxOkVYLuDyVy8SQUWCt6rOdO1xuwgbI77PMAoytUfGzEdujnMTtv0WhnAHtlTK/1cQ2q
15FHbVOO+Yqo1g+uSVjYQE/EH3j/qXtQCFk9OkvR9+CkvwYYbzWggRLfQc6uj3INlmlyy74YPyJQ
iykgzXdn09d6OHIJUbD/m0JH5IDb6rFOqf9lMXmSDx9HUfZayUxshWLluErUr+jXxD6k+E7UFHl2
ad2Uql9QVa777tcOEu17/0XQvpa14s2Uyywx3fqmNks44nL2FRbVS9pU2a9NWKj1LscThGRB2H+4
xrHrn2esIL8YvdY6eNzAcrxUo2zgC4mz8dA5Dv1fKTMEOe8cWQ2gPhWtym3Yz010kzKSF519kuV2
9Kv62r+jrEduvhBRympG9ejd9hF7cLXMSEYrUoTXPb6YswUPesjgPJcjBggK5HYaNm43jnFNwmDY
r3dXPe8v42zTRJHRW7L4llVRcvb9q2rb63Ccg7kD4Mkvlb+CLwDblYpm1inv9oL3pFeEJL2zgH1N
EqqKRx9ZOFraAHNkKY1yON7l9Jy2ZXzge6qY+I13sfS+qQktNPU+oLavCyvV4xpp8rIV3tv/x+3X
slWN7slgPxaJ6CLNRS4xHkP/VW7r0pENfBu8teDqFm/MYxirXtC7XHP97Wt3OjBDQ3Z5MIySq3Ka
gqVxLesE0uhbHlYmceRWgdtczWxMkbBtFq7rJMursGLMB5b+Rl61bN3YlNklbxSzNhZR4IqdabZI
V/Xa5YY8iA2a6IzIbHDyWwlGJcV92MwGOHOvfYsKMTH8/R3si32YfTiPNqi5lVu4Nl1UTEMO5cau
TMlQ3HRUEklU+KdkPSNWi/ODGQuVu7c6TrOeqc7GadjIbNj0Jl1v96vbdNlOyqCeAUc3D7jreht9
NGjN9y2pTvr9BeUw4WEcBJt8BeBbeO6hTw68KQi8W/V7YY9avVrN7xfE91/nrdoy7P1nCGI+9ve/
UAM6ZvmdQEnuREFzx65E0Pi8hgrQX677mVy6tloEHPdYuhUzj0yIBv1/ALLkwmqLfp/cUJEUZu6U
GDgOfFQUcUvdqNZlTFeq6SL4d6Z9UFLm1GaxrGyWVmXlBWIwRktPOonDHgs8sNqGVhIUBTXV/dAp
UQw6Eg0N+eVMY2gzeVGhZwOOANMzvNdODWGsTRPdUNxrM1Nj0VA5vHZicscO/iAXBZWM+/vKgcc4
+gFCTOSZvrW+dTTZc4tBZtCZxsgche9NXBVns1Sm6Wk4LTSw1nIpk9c4AzBP/4hAGrbxQi8p+qWJ
aqX/LcRcRDGqQcfMmszYISuM0dNk5Up3JkcXjYd0anyZ6nAUEFTOQcJu3Yc7S5i7hZ+pF29jW26A
zcXZ3Gtdyu/cOqH5/nQMc/z9ab8MiYrOySPkP30E0L+wZQpvlpsH9hxZD6pPFiS8jdfirknYSZgf
9o6rueFF4g56IAHzo1/n6lct/k7KavjLfwixvmNnMKMsHgDqx6E//2oJ5jHNVncxhkYl60nYGvUQ
YKoo+mYDqdKTTa1W4xXFHhlcWs9iFFM6hUOsspY9omkHIIcfdW0QuOEROZCjiZBpzwsnuk5Td90N
0Cf8xvK72rEPeFV9qahIEDAsQAIHkjpTgBRieQOV+QMexLOvA3jYCeJP8TwdQ/kreAgx2BUFwCaR
Nw37L4nWMteHijzc0+CHJH2iDDlqszCblrrH8ZUCGFk3IjkiXGPk8zKON7eznsdTCMtiOJt/FOlL
yvK3ErZ+iWlIIpgBbBb3HPhgtTwJCY9FgB8ROGBSfsDPg4HfFvOgBlRxgtoLGDbDX60j/SoRGEoL
LlP68+E49qBn3zfBt+FMVQxyi6IcEeNiI6V9aI8An2ypCzR3WDN2QOCAePlXUL1cc4WTJQNyXWwQ
FmF4BmK66lQK3xZObRXyNmWQ9SMt9bFtLYFmGIHbOFint27AkAe48zEVkkdQZ6GGMr4b1cef6OAT
Z2tZCUieDaHcxnngaXo5nD2g38CDtSSAxFhlKnR/h8c37jFdA3V4NGIgaLgvy87Yg2tWe0lHitzj
ppKDIi89Q3GsxB90CN7AUENPYPq1iedhXana3p8bYlNPGTBy/UhANPWakMKzmMyAcNHu7xR+8KNm
8TNT0oB507sI3wSgtvBaEa+mHVv9IBGhf8gKImkFYRS0UpfRAhdOd+UGxzABao+4LDTsh3s7SEVy
EvGYIffdX5qHtH1kpkMu7/IZwRmI2Ni7zCvbe1AilTNh5oXSIB5wKAyVBlQK2eKAsusQwl1q46h5
dguNOy7/spDTZuVFZIphRUJLvNWvwMHFEATPJ3WtSISpUEqKKSdlrJBS57K11K2s8Bggp6PadgX7
CuwJ9eVdEctc/rv6C1LwO21BQrhP5/TNUZ+UC+tfiAH13eFkCzh2SNkz46nrA7GAYIy3fv1B0Rzv
1avLn/ckK/pgbaSkkpgvhvbZMZeOAZiCbi4gaxFfpgZjGWOMH0JkFYsiC2EUuHactjomiEPj6PMU
P7Arw1zX+8QX/FGy6GZtnRnGsK/oPFCvJ9lgCS4OvlGmqZQJled3R4VEZYNV+PAxseVzPlxYiEd+
LenKsEslF+5cYH5jg88pclJGO5ymQuNfTp0SHo221Q+xkgZfHaZ3jvHFxaJPE7RluiVsi18xJ0iQ
LqmKvSPOBZ1tFRDgaJiyO5GI5aIlRydqM/P4CWkiqIYo3bvtAH2Qh/o9zTYoe7YLhs9Y/TqOCzGk
nY5wzm+JhRP8OMVrZ3MC8/RERQZht6oCIKXxKsHERrQjkse1txeHv5VlT8481ZSFNvDnr9QAjfGJ
Q8S5+PQr3jF6Z0Gj348PAkzgc2pbwzbO+QrSJn0eYHQAEzm5VHy7i4TaXdfbvWynkEJsxljGda7H
FkSOXCrLediofGAY4ph1RSyJZDaj4nCQRfIAPsfAmasvSp6GCua4Yy4uJpJRIYvlEsqGE8pcw00h
xBKR4ffCOhbtT0UaoJlQRIO+ROxz7XMw6P+f5XCky+ndwrdGYVqowkdCEb0/RzwKFaREYm4RdIXe
6QxM0eBrLhROo+x/UGY5MYW/e7l4a0S695X5s8UqEfEGVCytf9+HxvWKBVkUtJqS9R7F/mgJjbli
hB/dSzhDl9gMwSDlfs3CVB2XHW+tmsPXGp5AiVWTfWPFGRxHCxIyyTKraR+EucYLyN8K1HetlqdG
iHLyf6jGbOKBpP91nQkG4CU5ndwtVxT7NY731aSqFqNpHQ2Mi0OjZZK8kaFb72vTkQcNrEVc16KJ
bkZqrdt/ZgHE1CQQ7T/oovOIZl5yIuP35mDwOysddew6NOHGf3Ly9baFaXv5v5lVgXV+9tAyesvS
Hi4bBNcXX+E9PkNn2CNdobCP36V3aaCZGl2x0+82oEmJlqyE8hC7YUG3pvKe83Ei5Hbe3AdJEl+j
TwRP6gsjG/1dtHxZPUoEjK/QCG5u4x7Ig3nyNvEZXkiZq9Pd4SvtuZlrku3Log9ybtNd9B3o+xxT
eaTHiLBbL6gTkYx6OOn2+gsp6zyW5k/GGOK755lzxiOm7SdIJAsNazrHX4nI2i7n1gjpQ25jVM/l
wAB8PDQ1Q9ewsb7n5+cwlCPvfSF6wb5nQgZ0/D7+zA+S0vYZhHVMxEWOuXoTe970y06Ck756yHQU
zI6vtc45r4aKH/V7bdzcPVzDGPlG5fU/JIw2Vh/e/namqw2n5UcSxWfmXOPVPfnXnP7vepOyoRKS
Posqoihj4qkSy5fVUJXzpZekDiu/xrzEAL63y66XZVemfx97AIl+/j/c86lOF+fY9byc/RXONGRr
W5hS6kLMgbRcJXgj7ITEicDwJM+xNMG9NdjEFK+daNiAFn5fXsmhGCKhRPtTT+Dorgk6Nl9X+npK
69+8MUdpavnoTsr7mbcL/vF83SpGBs/Ojsyk9sUomftiTtab/G8humP0iWAMFf/nUJdmNFgWPWnU
FLUBSVC115YlFo7vH4OVDSkev5NrS1K4VTjOkIHvAEdgrchKVOQysc5pqUf0S2Z0N1Ku0N1A1Ybd
zjmxuEE+4vRPAHYJrYNy3Q8bAqkiMKTwhheHCQLgmDUKcGH6+Y8c5EiyuSsXZWWU1Zn3XoVoMPwX
trwJCS5V01JnMuNnHGAc4WVpA2ZhbrQdG+s1ApcN2NJxPEkAJbjmHCQ7RnSe13MVr+H4HiabTjKC
jefAx8xK3qA9p2gSoyYhyqmYwkBdaSBt28J2SLW8zBRoPn4W9zM13Jnf3cvVbcYjIk6MHQFN1Aey
vzP76lbNpc5fEslOmqZESQFMfS2T/j8Ns/qRlMXblKqNSkd7GdqNFINmLUlw8xgTytTHKSCh6Bn0
2M0TEBu2MG9KAafL1CEzVj+usOaRMO9yuZrYJMzjML/BsFW1eOUdTfyvCc40JDC1fZek0CxNwB7M
Q6jV4uXnJV83cpEjg3tGsOaNJE81y7MdA8qpEnKkMT6yh+ICnK3t4TuKFM5mAF03/2zSvZbWxFd5
0skrvcuQ0i/WMgLB0gz1w4+AiVEBF8PIQMdBAHfgPQBIbKBOHn+HWUxiSm4usEckLVX1gNNMDBZ6
Wb44a/PPKGOlyz7QZ2bf4dILnvHvvKQDzPZOs3J4N8HyBNAvi7r5u52nhMuBGeK9JugEf6XftmdK
p/ynA4y5mzK6WH1Itf3lasBYuazUZMKadB5E/SqwYVA11oUGpzCN71UAnFuFihm468FJ2AQNLofx
LcQlQwQRDO5PG4VuYEOd+zjATvRG6xfMGW6xIjX94GI5HZ4GpRaUedeN+MWNh9SiP9S6W6VPiYzv
CTu4LT4Z/Fp2+yVSj/42Oyr7m/grpWiCIfP9qPlzlkk7MMYxVF4+gHvIYG4Rhcjn3Efao1d/xMih
hcxjnX7C8lYZktZv+KKyqD73HgfjwDRhQUhuaOO4RBPFrg8j2nf/7d2/ytHF2j+qFt7Igz1pOcbo
TGUIEYWRWFIoExVVzLOsSaUbCu3tTesu/rOCVkYVeaDREYGDf0WIWzjF7lIE9YH42FE4BhDEvmT3
3iQVqWG3sLnepCfwvPu5VRswanhzTMgfFsn9/BoBrhtKsdhgrIL4V7lWcqQd/YseBG+3ZggGRU1K
urOICMfpZHsd8fvYGKeFz92PgYwNrxM5PSzWO74WGo8UDKWplfUTQ6xTJNc4PJqZqHWkYlURLQZY
65/rq2rZjpRH8BVtPPnS9pivzvQe7dCC++1EL9o/kqlF3dvHcinvDwd1zNhq8JIXtO33CHwdapcM
bqGvT1dMYfIvr8mi7p1n5QYK9mfHThxVLD4ivK6JWY/ktFUw0sLusrr/tER8DC5ZMrelp3N3sru9
RHgO8jkJJAEl00+fSbqzk9qSP/j6rA0rENJ86aeM2I1o5GZt56YlufwR7wYSyTHJJiLntJ+iixa2
ntBEcCXRzf5x6/oteuSZI5kKU7LEKVxCBsA/PrBcubh9G4orVcCp6aGzsGYs8js5nCgeAux0lR6m
cD3ADHtev80bdEFZi2SL+T9RGQvpVWKbST4oxYSF20PrGv1qVdNv1TUVC7rL8yYicrCT/UbMvC/t
57v/hp7V6FmYZ3c4IW47bU0OwkP4g4+vZ/YL42q+Rm59htqYfQZVXiLjC5wICWnPkbndKwKhw140
ZtpR5H/vVCnEvBI1eVI5+c01rrKWVCWpRdWwwUTqS3iQtl07tf9l5zWUqG4qOsiXsKpOYWIdBnnG
PVVA78eJRDC0yHiA5VG+UY+35PdSOMGu9MovBjCBL1NXCc8lgx26FjHBqOP0HHa23IHnmB/11+6v
cjYnMuNsKrSky6T3uy8dPi0750RwZnn0PGoZu0RV6vekOz3scl1uf8oI6MyT1apWlZexeazwfhR9
cXYhQz11rcH1PRJVPjWHeEt3gzYw0WwgP5HIGYToztzPgPdQL1zsOfMXWid5lS8khbTISQRvuh1Z
0MiGqMpR5Dib7J+Dnyv0zb/ledFbopXUC+jZU0IG75HHUqqQg02598p9inYn04Mi9IiVOJIlS3oD
b773qFhFJL675Yss2O3u00uNpI/o8ZVorhKWv90ZB7jVtnLy9vLUFJDJg6pt611eietIuBl0Iv1p
jryvZ5HbFDFIryHusKlvO6vbS3jaBXbSy3LhJaA2gu/bAfyBKXaiDAJK/nj9ikE0LTsfqPAao/Of
jTqKRbRAFBn1S9Zn4y6ck2r6Q6Kbqlsd4CPvnec6TMCUXhrx6TSd+f97u382TIAouoSv1X9IW1jP
FZcb7nhQZyBrTjgha2a1ybg73+1ZVgs9f3QlaraoOuJLesLi+Q5qGSgz9/X+Y+dpNgYlfv9LhiIT
9H8YWTwVjYrjTmZ5xcQPGHktKarAt4zWw2G4EpnE9poetbhY/0qu6kAjTNnDN7L7kTVX06ym7lre
r+K9e+lfzXtI+jO9zhaoc88A02FLgfDYzLDoiExFYOTW0pVIBtWL0e9RKB8m+B9vcIkTXuY4jdH+
SKKUH9YbuuZyDSD2ZIv5Jy/6lJISPVVrqvvLXvhx2WmR9X6SQzBxvGI6UWz2Qpv3MEd+ay6FzQpS
8RrbHyhA2wS4p/t2OUJwL0cc8f/ewW1QBSavNGAE9k2F5NbNI5HqIHaTlV/743sCEosJT39QacSd
A3ytZNcY148v9Jw342hX3i2ipJy2ER0fA/jV4SZf5vgyPSW9aEGyDyUpd5IFXOMFK85VrwNadUt7
HDIhybnAZNRMf1i6qteUJ1Do5PVFsSJrR02LIIkk9CyeIfQr3PC4Re3Gc4UrpM6a7UX2elFJcnvX
5Y6WIBQYvnJwmMLb+blB9ity/XWfpuliuUYNyZv5WqyD8LuAKkEFpjLzckyg5ldB3XxjBmY3HYeJ
KsRpzBmppOWbzA319+XU9jtCYdE1LvJzVg57CObDwkyKGiNOjCimVQTO8MyWuetXRJbuVusGdtUm
T0MbLBHrxILhKjB8DRObLVqzaM9hJ8FOPMSsgM5KL2St6Sfri3matLRfQVhzz78PTHE47dOn5ozp
lrUjF6QsjvMCckY2BNMEVMpjspmRzUydTqSFzsIlieZLVzzl92Y2vNbOZrZeAcRJM0CcxM+igg/G
87f38eHRdeOLY+NNhWGseXimfE6aBJa/LXXiBxVONOTo+tPsVLKBjqZ0MqexraQzXug6KkNHNqFi
qQJqhhYV5VgnukrAYdnCrKjtOPpOcT/XmX6TQjBkLPsDq+r+We1dzqYhwti6S5h5CQtqAVIzxEzt
PF/K98BOikQH2hmOUfzzX/HFIWjMb3dMjROoMuzlBKp1HgJoyMNkp1mKryUxiuzuJ/W5X7fwZKd+
5UhyMk4E68+Qb0Py6UCy54hFxZw4JQT0B01tmV8tx/AvtNoHmhgkY5tHF0QQscNptNzm+oN4mRCy
KDkVUlEmfBAFPFN5ryR6Vg/MYv2dwf0uNDesxKrDackBAwpzGfpX2WDBxgxQn4vvkSSjJLoGDESO
Ej/CyRLHj9f9MHMdYLPVj+CsGhyTjEBKoLYqXZ7SdMVNpGt5BADFo4Y1sgPLwOYmBNNvJwAOdiCN
+NjdSsumX5dlU8TInfK/GkZiNMsptI+iEDYtpLs8uc+w0Jdc8IC771Uh3DWH55PWzRzMuL7pS4bI
1S3rjzAmfWF9b7e3xC7n3IwuvRG4aEj8dewGF3TWgFGu6+lW+DNbXHd2H8asmD7mdllamTVDViOp
PHzxkv0dEtrFmeoHbrHiEKMn85i1JyL5O+fa7h7HtmS0lA+lx4XeP87WIUY5fRRDrNUbvEDnfMbI
RHAVTRIa+nS4MpoWP25qenneAqZsGliHJ1nl/fZsoF7/7s+Ma5aOVwxOv3ZKLiWz0/GOuxXYbGgx
WrOVIBq1A3HrhgeP1+rjmH58xYtq3QOUyNfQggl/7oqHFRD4Y8edpt8DttZJ9AL5g3j2dYtDo19p
j/oaeht1m2S9Jy+EE2xBvlUidoYKXo5dTv1ZPNEsNsVVZNwynuQNaVI7xpzGJlf/l9MKiIS0bFd/
PaEt+quWx4PInPjA1yC9K90XZxb/g8b5/r0ZcCasWwPwRnz0xz9geBLRc5ynOEifLQhrNIXtRjfZ
yArLum9CdcvN4BxILSoo2ySFTrFnxTEGBzOMshjFHT4nzathsoX2MeUWk3F4zDIQtX0ZLE3vgZvs
jAdxHu2bdlOmWVfOqMCdvpF8bvOOhf0s6MUWZYINd+HLDaMSUeSwujwK9ld98VaI14xk/h23eqOW
hdJX3gePvAMvMwevMQL+h7VnkXAXor6F0WR6Q/bZjYFBCr5WRo0eQUgA4LR/O7FX6VLhXzc2X31z
DYiOkRZhb1kCxMx3RD2XgCa31v1Qxm926Lhx+eS/93/Og3DHiKYxHjwqugplR6ZImUug2KYFx6ar
OLjEL+f51fHHkxBij57A/KD1+bsl5Cg1visRPuWnAFHvGKFMZfO4UyJHQabSz78suE4D354GpZW9
kIJY2ezcFG6uc0NCfjLBdyQETCj5UUpC1j4Ep+9eI7rvEdcEvE8pWRaPNF/Ri7Y39aI2hZCpnZbx
hg9W1S73LgZ1eQUhfiGLVifeRs2nsP75MizpQG+Puw2Fnj5UWBbsVAZhvZEesbnoVrvmB/Nn7iSg
2RYyO9SMkNFt15VwfTMisj155nGLK+QTYuuEDAJ70d499itd+UuSX/9K4VNMYMRmERPPUyjixsQY
ja6vpuufDbFIvaFOYzhBsoQPL2zIJC2tBeSLvTkekTX4na/OOzom2vs9e0v2arrhuspGef5AppLW
p9r5tHS+IGBAw9ITJPhHiNtUqmfPEJ/f18bEmlXhnj7ESG0tUsFPPGBv1hqvu38ztajsLzPjxnqG
nKOl5XtqzS5N3hpRUdM48v56B1gIlQDfeQ/hmvAuHg56LyrTZ0SPIMGQDU90pCGVWJOdcXIaeKIe
JRuhJbctxbR+IogodDnhKSpa9eKaIafIrjNj3nTCAYg9qBhSVIMz4as/4sg/aKoiOPwE/2w3djLp
BmE8TqcVNhsp6VT1Sd+4wNTPuwPgkrGSj4RAmw9xvjpAp0j9qutYAAxyB+9/x3dCkNG8Y5w/VxXc
DbZ7P5I2zNG8wgiBV7lgUOJ8E2hKkItCFsVoYrFfVRxG4G60xev4Cjo4RaBhsSnEBxdRZ2PcuGZI
OeQjtlbo1h9qJMACPg03F/eAwW0IlYD3WJE07Agb4OtSosxaux2Yp4IQiRnWtsv6blyrPPckIl8Z
/YQosWUcrO85eR+dWUhONd3ewR9tPqKAPJe82OVCMYuvq+DQv4v4AM07Ltm1QF4eY9d31MPek1z8
vnClchjBhII+xaJ1talyedFJcbNs97/zIMBIAceAO0KSSZaVxy4FYwJUqGScjGVUxcmqnFKsdtWa
trmeyfP3pEeZEaQgO6a3UMf9tOjmHH+d8xPmrpVhrHIBJJsFLasyIBCsZ40FNhujUhfVKzj6yfXW
UQoUCA9+lG4ajlkTnrTWnSk5GwvSmQuQGyJdfroluKhvt94BbKtTB8zZwBFL7MI06LhcnHQ2OlP6
oqunExErqVNm5WoBnZLTTm3GRwF79XC7ef/XT1vdaGL1xuOjfghzBxVeglg3csa/r1LLYYSQqQYO
P07MnaZk1awZUgNR1OvWJHhyJhvbC8e4zU/kljzNyhhzC2O8pPJvf9/xMtoxCczLk7+MPI9Keicr
zbQ1OvecEmhIfFBgYJZh9xS95vIj1Wm1haXsgZuMKLYE549zA/wU8ObY6p549upB+jjo9bA6n0kZ
6WG0hlkRRJQuEHJW8ODsacM6c94L37cf4b4dAETepdeTgjGyFUY2dZtFpm11nC9wwGwVHZwsBMr+
71Lb6zQk6wv+t3IlpcGnDp203FVud5H9egNW1Fzq5vjyRBgoNpAwvwq6d3hwJGw5l/iXY7mc/buC
m36yDJ/QkDeVaGYNKQGSmDQLRNMXMotFTcPtLLaxP2lOO65uBuIuyGIITrYkGh2aKHzuV2ruDFVW
9ydueubWPUmImvj/Itg4mXmy34Hn5BWBXOqjNrtEDasGe4vHR2C5OnvD/Fp+7TVKYnoBpr7tXw6K
t/RHrN9BOZccgxJjgVK1vUcttw5uT0Nslq/n3uND4mdkAFv1J7Y2usA+Yvb5CskBFVdD7Mm1dBRy
AUXfo4oVfF2fE9MMdutvzSEizMihbb90bDYezjIR4/iOnpsaeObPF/h0g2CZg/ZiPbRk+TmoIkE2
7SjdWWFx2OKnxwWrvbsrpLRAKkBkWWhPHJk8BrX73tYyLE2hblGLF9e+68NF+ySVusF3MvPxy2o/
Aui6keXLo8wXdDzPd5WqhoUSr9y8mI/hZRRWJDV5BApF4XNtEhlzoGtpIZSI8Ty/Zm5hJJiykECb
hf3CKemtlk/Q2vAgI/Gk6ITypsia9Dwf0zlKKl6F8UrArisVDEP1S+Sd4Eq8yf2dZgYxdo+n0Rf3
9u2DfxljrGCQnQGqDVXSv5jUkiFkLg1rpv7VUAqhvB/S7sDlZ6HTjP7rmwOlSa17zB2yqAcm9FID
LZ+i8GambizLNaOvmv7/nW4oUL5AHX96ev6FJk4ETGjUGhvWXLuz/ZJbONsq3D32Ng4fbj6QWwPW
5Nvj7Cew7pwIakrk6Ben68mWMlbBx7kgzVoCxcvzuGPfSjr1TTsFAcALDtMpiOEi+zS4NLWjDt2o
sQ6fbYcqNUUKXc+pFL/nnQ/e5Pz+6/EZEnsTobm1yn0Uj7f9kf2BtTxQ2/WajOvMSQeg5BlGdxqo
VzMlkQ1cZTfWaJ4sXGBe3SVArCUibERUw/BEREapaelWxYfUxZ0iB1fVc0z0qgUdwRhFK0yHJb5u
vHsIEME1K6iV6zOY1hEW+9wLD1qyrhq81eRufbGi8x/iRK+3amtUpPqZtmGTHmc9v5kfWTqzijX1
0mlfmW4j7SnKb4UM55UxslcEhq6om4Bk1vIIVQUkwWQwWEQ3htzb68aYaPcp4NeTxKYBUFj6UKrT
BHArwC9SRJTCaqA7ei/Jd27NoZtrdDLovOPb4kvcMgcyxa2SiX270zSofOJiiu4cTZODC9hYs+dq
FZM8JPR7MqKCCpdndMQwkGlPI25ht4Ah6QBgAvzdsER5uneXtXLdUCicf98rVNRJc0pDC970q8iO
BCM1vpwExoE7ubHgsMPAm8z6UbvIGLlY/ZzrHa7emvJbyJZZ3cqVuPyOZNT5GLkapkKmVfGMTTy0
YZXq4p9U4Y5SsTc+faG9PPCPYGu2SlAqMyDq+Zj3ehGtm8i6pzDuig/lhIkb5fHteI3gFh4Lji78
N2dJWFppGuYVh1A9+QEqcdW7Jz+67B5FsHZ/vRXGSvVo2L1LLx4SOENSmGzU55jQShx4JmGxYbvI
MFTDzt8w14ieTp8ZRBrvi1JYuzBoT4ldXb6sf5tHCZPE/PeNFbIfJ9eowFK3U71xT7Mk8Z/+6YvM
zqqXVB9DXrRK7MpxUMyX5zhZ+bqMjOFp70ZLuKf6D1HtTDE8FEf8jzA0PDbRcNWD7vSPqRbd1dAi
6ybcld/asnHkgd3dE2TWqlWX2S2OeiWB60Z76a9DW0gQDopJoDsH//AgmvekmUZJfRxNPD+m62vD
rtAEP7CyuEpMxW+HhmVQHVL2AbpbaxX4bsapc4BjoLsUW6L6yIpPVzlRantVrYFeX/Q9rPHOf+jg
bzuy6PSjIVFAOxVLq7kQZAVWtlHXo0iL7K1FhrhqBaw5TaeYL7l3eofiYrj0mhBXf3NVgJpu4L/q
zGNENX/YLopa0VUaVz3VX5+q9A5mWTKjPk1QX4ocf4jbD3mcct6pVOpMSV/s7C4mJEwRqN6BaIj3
EW+bGkucEAElMiQZT1vD6n9EHlfEf+y4O6Z3KN7EN8IfDMUNfze0+cYw8dEjEcdO3r6P4Yy6OcAR
TZoXDxWA7VAie+HiguoXk9a4Nb4cJglQqtzgCCJJC/KeSABqCb7JAoAaKcWQOsR+DX/7BumiT8rW
/ZlGlSsKgxIc9cwUjBzmbpbUub0t8WUANXbols4S2u2nxW04INSjdBMQB2SXxxAS27xYDGWz3NB4
IfxeFgD/dWG9N6kc9aoAGLiqFkc+eyxMuqGY1/W2uWovxz1EI8gILBJjqJv5taeOcjjZm8/+2spz
Cw7AqUInR2R3gGMYbKbQsSqfWG8YUoQgM4e+ZMr+5ftlsyO7FeOs7iPus7/zRt4an+XNJxA/gpIY
WckccJKinixK5Sd6rT3RaBEeXqDRlyFsCjfQZY09B4IDMVUIf1My+tq4Eljezosz5ieVPrKM5/B6
ZLrKPh4S56zgE3R1ScO1z3W/lgYVs1s1OxoM/4V3MDO/Ogvdh1MQTmF8tK2Rrej2KtkVynwq2ikE
Otr0xx6FgNuUGKMEcxJbTuKcOGjJpyw5TlIleeH/y2SXIT2SPFXLGXAj6SLl23zwSjgoBm7IcZrV
7b1Bfq8yLO9QNEqON7Ewdtu6MEL/8vX/QTPjQxcVD/c1y3xuOJCxkcX4b8JEjZKHlu2XI/Vp4bPb
Hpq71MqHTn+iACekPEYOCSAzHBLrpp2c1/qTk9HNnZRgSH10SXCrGOOvBnDs4u19LE7gTSrCjZjs
UN/ffBPUKa+0kC9DFKK5YcSfYY+SvXrOt8Vn2gHjKCxGZCr4l/trQs11ZiJl94P3QleeirJ4c4kL
IEZwteXPKv9LpIjFYyjqUSJKIijXsTSHTTbMGuNkKYRVo2DiH2CL8QlTLJdmP9/uRLr9R+UGUsqD
mUec4igMPus8zU3rRLT18UZwrwvVSSrviQ8g5CGYsjKf0kieFlmQQJvPVq+suR5SwmAAWk20BqDg
FRUZrK3/nIGhauTdKZBq1/SuegL/LCreYB+oNT2eKmo40FnnXjdkKJms6tbnoLMnSMjUGckg0LiJ
fQ5xWNmHnKJU1GPWW/mdMCuuZOzfNpFjVBsiqqNNnLfygd3JrHFaWEaO4V7gRDHMTaJqQ8H/EQ5z
K5KAWciYDf7N3R8O/tftI8KacAj/tcMtIP5nprlqewQm56A4oXa0j6DKszIY1xJ08B4jCMcrmvcs
8X4MK2Y2Yj7THeqtcT/b1vj3UBD3TIZ+vpNQb1Jt8iiLBIEEjgMv3FU0WMtSGBNysKE5pmzsKyMj
PrQeK5+6xkUvuVq6400SEpldWS6FLmICZNpNqeFvY3/Kw9VJisHAD4eTJJh6vq13ILGEUeecreKZ
Rx/2iPyHw9paI7yAXkeYjxWOk/ZL8Oi5Zg6XK0xKZR+B0FUZVAa71ZMczmwUHQ/9YHl7wS75W8qN
TQn3VhK342qgJ5vktewwxVQqsR7dwX+Agn9X3WYHqIB+Btk6q2BL1kRQZyPQJvYuOAaiN4NNNIdO
i8CJyoLBTDZhBMjg+B8Oul+5l1eZWTJi2UJAto+qVYB8UWLdgFJT9bFAwFZoUpFTKjpeTFSkUqzB
p5UOmaXqNOU+nMHVtIp5BMDjHXeqycclYqwjE1lp2c55JITTQ+RCPFsmuMD8o20srOXBtzsx3ZuE
lIa4ve7fSl7X4s5f3qYLT721b86z+7/d2S/rmfiRCQ6C6e0OC8olQIyk+xDaa63Mlq66/1i9O5kD
0kQiZIltxKANi6QJnjbvrm0kHceYwQJgKRp+fP5q3kUCCu237U1oXJxEMwEIRtZz9e+eb9TKpKNb
N8JUE7jTOALBw7722Ce1BirSg4/f5SPassNFDNic6igdi0NbHxJrsM2tB5kCUGRPfOyGjuGn6On4
gqEjGC6wIYibGg0Miy8hG8twbMhuGmmkMK3QwjuXfyCIjkljHfQXFsFnmZsng+br863ABXX/v6j3
Q5ph+RVOKbUtEs2CUtNFeyGSJGVukpWK6q8xtVFAW/oiyBysIwUbx7IoM6ltLqgwH2LCxSXLUV5b
trfJ+WS4FD5x6fyPkqvRb7v8Lyt4Rwmw3Z1IsrxX2xF5pvZfeILlh2DF9PlcubIxafIJ6TadXGkp
UYdOY4H6EzhYyWamCj8gAAl0yBMyqmbYkQB0GuUThoCbWPeMban0SpWsSAi47hsin38OdzLkf4Te
32Vcyqe945B7guEoj7TA3rcsD2z7THKuVxQegPCqh3+Xho3HfLsVVzGSQNEvGylpQK2KF7bUJyXx
XJkUomOGjW/sWoLYH18nWNNSUp8DEVq+kZFZj0cJCUPXROUqtZDMdPr9u+nLZ4dFEMyjCW5A7aMR
K8mJ/7zK04mux2oMMpPaO6FdjJk8xvP+L/7S04hL1ZOLjQggJd1MCh8LrMcetUD5fBZEt/Np3FiI
Ujs65lXQkgMWe6wSXXryk2sLieSge1SKUW0pUHVY7hC2HkyX5zbuaneCJnM3Xqb+fUVI3uOFlYlr
qA6yLgCDMpQKVjTrpFGqLHlbX/sPHLwTbbblYFXGhDlzQ6P0YP6P8boMag5X38cD5aGBDEclQZsm
V2KKjH8r/L9FczZJQ6vUc2RQJIi/WayJFfWGuWWz8xZBrpIJRs0YXTpkXwKP569gEHcv/AuGh2FN
wUruBeI9w7B5KAVZ2IbkU5+YWuAy9RJ6QDcYLDc/WwTKojADCVURf8GobYmJ/d7XAIiZRhwfLRE+
5snzu+Ks8b5xK2+qAaH8R5n/ZdnKBq+f3dwVtQYqZu7T45zmtib0FrlVaDP1oA2TaPvGUpHQVFxo
hPz8YJ9Fpyn72wLOOjl/48gls2Yby0H6/O0DzUMr3Ckz4T2qYv7V97hEs1owzosJnh2goVqMTANY
F3MjRWlgP16g4aL+ZWHApLRffMJQjcp9xwwnY1ViIL2yJuHIyp+xfFbH+ZKxCN9ioDWshMnunkZY
muZjtxc83f8zzfjIsLf/HVYv5eCCD5e1w+iupMEgrRqF8qRoukq/UJXaC8pCv/9brPoaXlvFOZDI
shkDyEWu0Crje8L8W/gNlrsZkHZfJMn/lBLygmoH8BHsiKxbi1NXYnce0vkK7CqiQQ5Hyf0wNSQQ
CQp5IX2BAHL7fLoqXUDT7qFjcn6AUmolUcllbJgiUfJL2tZf1XELMYCaia+mwKN/2OB92jAIkwjd
UXnQVtFPTDKhuqR8TUAaCPe7KZxKRpuaKWcVoivgS0gcqhlCRd2nfb46sqHriqOeckp2z6GrVwhL
MlIrLodKWjIO0HkYBopEoopJ296n84RJ1mHVapm6JVexzcKvyhoroUgk+R8fqw+Uwm5xXKXQ8+6d
XAGzkd3RFfyvoMedPobDBzuEDK2U+oTdKzduZ1kB+ot5137Qlnume1JbM42wP6o2f4pkI0A4CI9Q
2ScP3RkqmO4rMkSZGS/QaXm3s9l5aNsMHBJNFmo5SZ2O3VFOd7NKzb8dz38tcp4yfUiXy6L+J/48
l8NjtRsCJOfqhIeEmScpfS33xagysZ6HXD3ZfWhZSNezuXm0by4qHM8V6GuolspBw+aCAtb48mQI
xOtdfZsBoMz2PR8wuiv2ricptWDlif9RuIKBcik17ZPicruKoVz9BgEl15X2koCzbwq7CTJnbJks
4LPKyR8x5Xe66LYq2xQ6NpzE03I5M497AxrqoN7RRqRhPRj2qZa3CrKoQFWQEoP7Ylv9XwMcXq0S
mW8sBY6IBXlPDitgtwe03DZdRyA2Rr6WyplI6CIBSVNmOyIV/bwdxlJs2mP/sxtFo1EGiDWURzW6
Wj7fndn43cymUdLBYDxwyULpAKAYgt30V7ecGml3zLy8OMVdR9YMsaA2gPlJ6kF5nVp2miBIIF5n
mSVLnakKYbBEs/L+jbCI7fkayTkfJZrCHn6+uYBOZOcVUpuV1GbG94uwv7Fi1VExdMP3cRVOmDyv
dh2AVBiI8HuBP93LAJWGAvsN/X1SbHDLa/1CBT7Oelte6LHGfAqIz3vuLzKI+Rlfw3vrkVe4HfGo
1Ss0X0n58D1e2rkxue2XiolSw9pc65CkkSxqiYPLA33m9m+PifKZDKpl0MjHfFdJF1uvjkNnuc1w
mFjQYr7+SoSjkJWkm90HiCKgzrQCW+9z0zLC3a7d6LbxoQUkd4846FPjbz/yOxtON6wABNT2gzXD
O3CabJ6QY4mwMzf7vXN8X+onxi9PgAAVsxoQCoUrDqgTdgyyNMq9MqxDXaVs0LVwBAt4pwq1s303
webH3PmK3ylIqRFThoQ95sXdK5L/cL1agOh2DVi9TcF5hOrq0gX76tpACEiZIqsq6yL+fy38maEq
OMMZoFun9g/a7qm+Vy9TVL7dGjxYcvMfztEEhf3kmvXZ4Uat+VxKxD3qkS6fRf/Fi8iu56Qy8TNj
s/F5iyWixol5uXHvKU4NtGs6I9bJTYjFjiU1vAF+6mnbONzUkiuyFkYji0Lt3qIRW2V8qjhIOQRc
l6rgTaSYqAK/PvytnphRzzBx7Czp+N+Khyh8mSDg363QNHEu+BHgrkvUEF4EYv3KHnA782nlue8x
iOzJ3Nyl6zLRir/XgqoLQQhCC214Ckc/siHWmFZpzEfzDfRX5G+mmqqiwPWcHgqjjfb3vRx1ejK2
iXdydKH703BH4mqHRrnTljN2n+TScG0mF/f0dvM3pepWkHR91AzhE3JQh8zXgU4PfLybdAEVBLrV
2yky9AD0bP1E77VvOh048QGXwujXqODjLifzfc1tTjwQumOW6vlYg07cKWqIKFGrS20h9XsRQmCC
hZiSiIfkIC7XB2cJewz+DbjqyAYSAueHzydczyErF3pDno8raVwKGum/WOHzWTwQ/JoO+5Sqb2f0
FPytHGwQAu35QOgqARvVcBtXL0yhdL0mgnPXoX82rDxOR6UJcHX3lRXTlWMxbjENHWeXBy1Zo9eG
YzDZchqtqR6B+90w4NpmqD4fpQ/3SqYLyxKVGr5BbEryzEwgzJsYHVA0ej6KpMjyqXVERRr7BitM
w9c0FRAN+2jFWW7g8AAZ7XzdBfl0H1u5LZSnxmudXR66uiC/u2ILsjYURFgz8cZMqOfHWJFaCuiC
oXP5kWeMOGPnKror5Fu8AYpI7Ic4w6TvQ426RdO1fmIB5oDF1TJQW6W83ZpByyjaqD/FeLn6QOlV
kUBAx4m6/Az3r02eRHmy/0m/+tqp+yws+VxEClsdQKbUj/4ENY6PBIc/vdUJIqG+98OkFV/ogXgT
TgUM/QfBASJSS0xbx534Ss9tHqrqxOZLYUqOFTdoLPd9hAfFgnUT0xr7AcerMJ01BXqKwrFt2uHZ
5+5h5TPaK+Upp2jvvzAAVQXNpn0mMESi/zYLl4uJgQ1cyn+rZZf+MYqN7+TTV1atYRGWqI/4o0Bl
OH8wkjqm3zFw1+F+FxopHg7sHy06LzYgcG8DqvLZHmpw42NJ4OasU/GEGHqXVbOj8IbL0aVCfcjy
nHEdwU2GxqavAGKTw4P8bE0JfZkmzeQRU6VLgCBkU8SDmRj+eHABI7KraA21MdG0tQ3jWxPy2ytT
btGiCvh2JsQEkLZXMQYTCxwEOQgS7M4huuyInNcDlFPI2kztTnhOkAYnHQ+FA5Au2/kcnccKqjer
y8qXd85YXUl939m2+U59/ITfPsBsRxJLnj6hbJ8c+EXeeGMnknA/2WD4yvnpN8pkDh5zRh8h7gvh
yi1p6EQA3jwqMLSuFe3yRMAdz5aRRUlDuNR0Xu8HwISB+WMbFO8LlJP+wFLAA8FDcORHRhhkhaG8
brht5RRQhYVcA85qbj41SYoGCb7eemNi0JtjeTDTygOaFBR1qGn7zlkl0QoGRQCcIC8jBPjVL5MK
O7Os4suzBOcha7HDjoXY0mqQYsd//cB8sEKUJCT6VHWLT/qylCmJTozsUg047obTGRbmX/239k8F
4X4aeGCIJaFHVi9NQ76kQY96bNERaOWN7+ELjxO2/7hwT/QhV4USaeamMUqucVZpBezY9R8LOVdx
cNv0nEWyrZfwDDUVkmZtN8nQfpRMtcLVBSErLuVlanTCwiSLiEMErSpW/dwxF/qXXQY8YStBS5lN
oozmEOB5ZTSEO105dim/MAY/U4ELaa3du4m1F18qGRwG/6J+BWX+xe046LwR3ieiMaZNUH/umju5
tz4Iluhva8CraisSEFnCqVKYcO2Fp5Wif7VED2fh7s6IemdOAEJ/TsgC7DaVv0iRiTUpYtldsjnz
CC+/Pn/sSue9rlynvMNnX1DH3d6FF2TCSMPqWfdcpsFANKwLDGOSzsE350KWN9eUvCt2P0w7zBvp
e8TSl4NRQDGfPCqMfC3iQCL7zLhWlYU3bIm0RnpxuiiIxVI39jLEOfF5MC31enAw0KWkde0BQjpn
nplXVduWBpzqlDQ0nhYmEjKCLrCvuB9SaKHbIHd7qxjAMtDb+gfUVTh9Do7We8z1SGcD6QT2qq6S
gI5Au3tbwFrm9/VdOb92nOfJWLDaxrZYziPho/5Z7UoHtriJ090Qw1XUgvv1q2IK0QY6+Jsb5jcx
ugdY7PkrXWuFdZK+dZlADfMYV/asUFCl5UCh0dL1p7qCNFx6ejxs8LbVEbIML+hVWvrHj8EucNej
I9XYzOgrUQvewMfglXmWW35HLaJOKHw5Y8zSGKXmFebBVfUUrK5r21BRbtCD4qgCZsUblJ0d6uTB
+jquGa9Y5YjBKQvY/SBcMBc27wPxG43Mhs7S/Wm+jXslxCjS5w5yyw/M4wpVvKMJ0TZDHarKkWz2
3+iwDLJWkJmONNJagCZCId1jsW96QOZQMVaiaajXuGw1uqWetGaGkCeNXRb9KqS7lODrtel62q/i
tj0NBurRr1HdpUARiQAy8yUNxr/tu9JZDqsfqe4A6ozjzLnQ9gwElR0gqUVekir2ngJAoWFZiycp
tmjVR59zv5uvTSiksBRAXOvzamzgKqPZK6g3PZ1fv3dBFgx1Spt1LmxdeP2EkBnUJhMmB4Mpa8KD
r/SYo+DAtySrWglTBPU65B6KUGeiHDd+XftwvoXqKQAzC5hfBcV2CfqvP+qKHF7lOChsLv5FDYwO
Fph8YTfe2mFycM/a27+mxjlet8bGIK3q78MsOD2zvZzcV5F8wYTTyiRwCsFij6qnNGHCphdr86g8
Nb3wS66uskLqrSy1adbmj983Q0/USdG3EqFmsUc7l/mrNwDQZSd6wc5gL95z0i4mGNPWvEVWrnxz
6DBY1mhb/tuCHGc7ukq4cArS2Lq0NQ39x3FfGsm8QARRR5+ZUP6s5ir8qHkOGrFeA0Y/54bk2ISt
VzGL5fG/4Hj9AL5eKuhi+dJ+00ktFZPTMekmpLB8g0VbgLAB36/2ZH2T/7y1Wez5kZMPttlX2JGp
rD47asK9Eb6ZcgxcVM2nySOLiCcLIao1E8nTt3/5ENFhYpRoFd999dQr5wHFOEAaYkVeF2pO6eSD
FNiEGTM7sc0g2quZruannxclf08agivdXrGOAdpl5fuwg0vuLrQEbA31GzIRlkBe6U2iamE8a3gI
/2mWdpqzfES8ox2Phes5HiZCxbk0k/3m/YiTz9++w728knonjzDyQEQcHw1VICtYbZC8W2mQ4Lyl
aqQj7GnQgqUGekSYRAP3WgASMoHhqQlHUfhHDg+ZchwbGnO5r+NdJ4Cxu1wRFmJjW7X+ZhrM4YxW
mVf7fIEzadWyoNSWniv+XQE2ZqN90v1zDE1Hy79yWJD8v3ddUtMgVoUvmTZz89W9rCjemqPqxYkk
a4bua7oT0elH3KvGmaNeHfVD/Lnaal5otUfzluZAk8IevVnKsmHTiqAa3xNSpDqs8eb3n2A+boa8
ROA9jBcoiO9O94beKiELX7QMN9QwpkLRH6FlDs0enQXuAsPdmdodIgaXDF3MNZN79+21a9gfoRr/
OrWMxK+58g1y0WyK6XMpqo4zvSN5PWhLJFw/xIc23okp9BaxDy9TF6+lEqXTGV+C8lq5KOsU1SnK
0hxQe1FjZk5SlslwY4fkg8y0CnsnAlzbRnv8rKQbP7eJiCy8pIZ1Y9yi1vTibZIIUYA9U4CTa1ww
P4ye3T2V+QxCTu1PUCZp0hF6ZNDA4zOav27NM372Af853AS4iIhqgtTlCvzNrDhaaCjtuvdJxUEn
RctULhQ8Rc4ceXFYWxALjFFWTldkdieBVOUGMxlIrEA0FnGVeV56UFyDlwnIyo2LtfNuplopzuTF
nx5aGVNmcoyWNsLIRk3V4jdleZ88QI7Ds950NrsGLfWPX9S2M4pw/dF0zYNFo1ZVn2A664DPLc/t
K+Bqv6dwbD6XXXUrbL4394FuP0iqHX9eAuAZqSvGZgKRffjrgPMoCqEUUO4wpsL4cHJ5DCkZc+ui
tU27S5aupi+7uTl/jB4lXOGcOurD4Rn3aSK41M51obWZ6FeJo0zmmC16CR2mc9FPnxi6apu+NHSI
TYAwgGZamTNd0uhSSqm6lfmJgqNClqVhNrY+HVwq+dMQK/Ih7KGsm6Y3fwhYwo663gYDWeIwGfPG
IMmbWlC4cNvtY3DXxnJSIvwU4sk/5H8sKS7icijLsq0l/QNt1bVeYsQVaiMbOI2zJBF9EKkO+9+o
aCqj5r5NRLPR0UuCI0Lxu2JnyMW//9MBzP6ZGb9TAxqZdxRVr93lJH6hqZcXHdSXncA7OD+XCpeU
W8hbRJmVeA0mUNqmNYbefhc44vTsQNAI4xxWCbRwv4lMWF25rd9gLiGlMevpQS1h1K79MONUR3Us
ujVzyw32NgshyUgKusk9vWshrnYBXBV6br4DE4ccTZXXoKv9PW5OxUR47U/v816McSvaaHEOU3sB
8uyEeczppQuTLMrlWKhlm++kOxEFal74xJea/pVPi4N6sXa2sz/qrgnVT5HncjPEZ/jsJAD8QD8Q
kWb4wYNhYsQOD7ZtQ2eZmu3iODjD+mB2OYW+/C3Ks+M+P7+PcbkKOms3BPa2h5BEWvVo836Jx0D1
C6OZ5O+iWHtP+1d4RgoJl4rWkNxjWdOR60EF+GOA0aVV6FSCR0PkNxrH6sW0GozUj0bUxybkGupm
Faqaec1t/W+ZVpvmIzlEE1CwrhL56W3N9Gu54szOPu9sQCABzttm8dQkUxLaHv6YzxfNeGHxD0ic
xWT1SWi5NCh9Nt7wllrBWiZfpvP6qh5F1DfFf6tQhpDCE8xPGaz3ZR1KCsgBr56sTNMg9M0OwmP4
qcwpE+9kVIkNSvZ7TVDh/wnpVsJ4J65R/OqHvf22fdhSBSFE6DSHTBH7fsQuZrGz6wO8RWJVOp7J
uOZdb+Wsy+Ow+RLVH7Iol79ULTBctHGQAR0TLLRmCu4OPEOk7g1pNDtWBWvtu396p2/9e/qUMqRf
B0t6brMI+nibKH2YCQqwm6qZNAh6Kr1hRDpMmaQabRvsUhb7Q3KnZ6ia1OKHT0Fzh1Q+aTOwlWon
JPjgBOQ0QqZl94q0DHZLyrvAb1pyQhxzzkjRSWcjHrmy4wkrZiUt6zhg0nZvDAczSxNulpguQTBv
DkZ3KBXHeIyE/zG9sbKDgsqp6DcRMjjyXprT+xfStWkHjXyCLjItAWukcMXLfd9cTWwPxWML+aco
/cXH5Fey45qTEqKXelMWd/R61SGxdziW5/upFYajj/MI4wbRL+6W0HziF/W9d0+GJv8Mzj5x10tW
1+Htp/QgXKue1MsBVB/tnHqEHghMur3KWaQLPeQKrjjMa4D5n0lBLwmTBxTEjTEnLLCfDarHD1Kp
fnIMErP0VLDM0SLpTJKuLhLykP+lkZLQVQnH6a23ocxRHSYU80w0LwjA3BH+tNaZ6czwxTVOe7Bw
vAap7LQ69XVqvsgVFipo8K+h2bBkGkpjzjQCNa4gG7I4hjRc83fRvs+guoeBVBJM6slhzGKc6MYk
Y1KvhW/8LBH2TUUUY0wtuuFjzanMpkpjwrbLa11OL+43YPf5ZNsJkWZnfXfDgCGnxE5ohQvIciB3
YjDV0mP+lhYz+/bO5rMrf8iYaD2v5Q+u/yWUPtd3NYakDBT6TA61FXRFBLFWuzZI9VBE7gZJf8b0
ZWVx8nb0H77AdOFp+8Y9ycDUyLG2fwe/hLa2fZjzmEPtL/oYejaqrXUmx2JUKYENniobCKlyhGiL
Cxke/dwEEBSCuDEmKiSStBQz98KiSKLcLLoFYYg5151doVnL9PwASnHLroIeuOul7510ZgEFUISe
ftcbs1yLBTtI3zsSyrtdGCN3p5Fi4M3tV5tljf2AMBauJBw6Sma3U+PTJ05f/dTOUE5RPojE7S7b
G5esb+OBKK8SavfWV6MZfSOeOVYsX1IzM8dw9O5MZTTRy0CH9yD5c0Uv9L0kpjj67Uzu/c/ERPyM
aWpO9+UR2UTPSANcfu79WI7p6pNUyY1jUxsPnLVtGx5zrtkpEeZG9LPMBrJWb6aJcD1zDtxfBdSd
mGc+C3nGrLtAt2+um++cXOICcv/rgPwor7fD/OYfslfS9EVjADboLGNDh7XXbV5O0dCmQDG4CK3E
/Sdex0TtNiTb+FYVtMxrHsg+RUoq1nccDjDpq0lxCyCqxBcULWJJeWWQpy7CbRD5Elo2zndet1gc
3P4WFch2q0jREHtbruHHOJxXqaew6MGcyqBVqgEci06wsX4dwFWgSvGjO3fRgonj/Df53VZsxu3q
P/BzkDn8TDR7NY9OA0vmkvTyN4JhjUqveUuPy0XO4J/g3c0yAR7lcr1t5dTCVivY3oiMZcskjRRx
odPcb9tu7v7vh9o0pOPZ6lyp0mMfSwdXnJtdQ0ECVDdDSlSQEpBAUhs27e3ICyPvESsh0SXC/BXu
EyL5t4blWJr725BL/Ur2mj0Lbc0/M7SxQp1H4QO5b/hm5gEgkUtV7sDGkx/QXij9o9kML+PFHSKV
u0AVhXRn6XFIvfd+DSwnLYUh00/WW3cViJON4q6TvNcOEFDYLvztjEEi48+R5BeoOXzpumi3IKMS
KMwW/QY2RRbYZNwUbODzRDspNhxMdw50YRg0iTs58doLhX/3Fu9KN0g65Wj8f1LtkIgDzMCBUdTy
DRksUX+EVqYKT4fRyMAkNCWLo8aSqr67nTke2rz/R0MO0DDurXEOREGk8T+mDIkBq7860zB6eCIe
v/YhAXuDqrNEugEbo2d/0uG6Vu2rLfYEWQpe+SQuFASedjatjwGQ96pLw2hroQxQtGOqTteIGfRK
paRJF4pwk/+eR5XRWL2b/KusR5wDZEAqs3g9Zl5oQ3Fwq6vGT+7RVoCHffJcKkfNuKBnj2RRpPRS
G7J7G7s0AxZA79QyRkPbvVNWIFoASOflc5nmzmYv5h0PxhA1lvWKGrlZ2T8KC8zTZKx9LLXdOcxI
QSIpBuB3lHQGVhdIYXfdwYIvUPUpJQbo+wXTBK7FC1mMLG4YmtqMBAf5YxVs/Q8/qLiFgJ381Uti
ejl5n80jxPmgKkZ+m2JCzftQyd3wdMqiHar/YOUGZjw4APwwh/JGSopoZLZ0gLHi46uOBc9foGYU
6b4wzpqtidiF8y0UgGfKeajwOwNWDTqRPqHQ1nOLde6nZb/Jbb9041qOG+PVv8yZ+LXHZnACK/QL
LQ3fnywGg28LqO8M9rJLU2fcpMO+SUx8v12nb92Bh/55quBbvW6I45MN+OFRZ8Hdgzh3x9x0Ll6n
biw02FnvTbZzk2+QixoqjPpeD0L4KjtidR/F6kADJQDPjTJ0DNkS4nPr7adC9zMisTRnULAAXKv0
7N/F/rnNouViWFavdgAjctpXA+IRFQKW+M9QbSHthpvRJ4neCbMUwUU0hHBkY5Boils/IN1YgjYU
joUQIcX7D4iyIX4QdWnhixWIMIYWZwJZhn8cfNYxX+WtBXIzwRYQ4iM5gHYq6MyfSDNuHzMRPH9d
WitXc2DvfxfWj5b9NRHMpruFDZjGI11rzmFugg0wwGJtNClVsXiqAA0irJc4PtDZb7yLGcoLozf0
+gYXKlfSIY+YX9cukv0YIncygek4ix78U35iTTGK2VdyhVGsH/o3JxomC4x4Ie6FYj2qhzffRgJS
EdUv3acFwgJIZDr08Y3lA3TWeA3uCkLmHGG5tiZbKXf62A1b2fya8uph7l9M8Gj0ztxazdanT/Wv
iBjfMgZthhBx8CRjYT0gy2l1NR8/l2JcaUruWlRF4iAGMSM4l4w1DhRhx4LNu/unmJ/H+KtZRIWn
VLvl7I7s1xgeYv1TjO4zB7G3nyIoWhfZ3hkGLzLHTFbOedahD4ulenPQVSIfnEgHEN6PiVnFKPm8
w8Fp4l+njp8Sf7qW7bizBIza0HUGmlAhBcLA13At1P30c30fHPNo86eltQsx6FjKmp+dRjNS92bk
YVbAPiDEVJW8e3jVr0sarNMaDVJhkAcuwbUpZeloaREdZ6fEe1GQt++FiHNDcd9tzOw7u6EUo/hS
2h7gR/DBtBGIu49lMPGaebvQlPCeSX6bJDZ2bS73OZHmW/+jOytm5wZNi9tJ23UItz5fF1YBcxSj
+AXnP6RA4dwpnoXhWIyxeFLoiwHPeoDhx6aAoB8f2YGFZSXNvP0DPlgFW+9GI7GR2e3YU6WkWw8H
X44ZXPKposmkpbActk1vC1SdPx+JYHtykmhulR3yfwGbwl8t8SWWpMSJ0Spr62aBxN24LV2W3pt+
w/JjKkKBw1/dPlwiUQ35CeG6QXtd5EpP7U/1nB0ICQxIM9A3dKobOCr1/CbUsHZ2pEq0+SD0x0YV
yFxxpn2wYY4J3h5A/Podasu9mZ+1+B7NmDtZwsYzzf2NTX5nqCtNhxp8FObGYdACIqfhDNlgmVbt
PsLU3jBkOYOX0ss+C8DeUkXVZE1Uzc8F5kTI77Bx+ThmcBcYJCzzLh6oPP4oYqA+QfhkmjA1V7XK
p51jwP9FBcV+zKOV/Mvwcv/rZN2VcH8HNzSCWxw8uE5QnvnOylQaGyPN2lD6JXRbXg23pCzFMEvN
2/kLmmYGoWpqAdY8O/9iewF4cU80j/q2INKL3pJTs+IX3p68MU5l6DhCASSY357F5Eg0WwlONu1Q
35eKLucVz8djojx19EPNEDBkXrQR5uuzY/J5vui0D3v2g1CmXDh90EslZdzyErRvIOVwZ5qccoW4
bx24xODoXvCbWmEdQwyEMdm2QzYJ0ZkdTlS8IR3xMemNChzvVGlc6ZKlQT3tsUq5BrrpbaAMwNUO
6wMPXKqd7e9UKedtyVqkkAjzxddDpKuLMt+TuQa6K0ijrDkoRb0V/qWQZ3oqQxLV649Z/iG72Z8T
dg2W949GTaXxea0aklqI5qoYu3oAf5U2NmPHYz2YDj19c1uDDvRAMD7xxYplyhKNUeWBnK3hp5R8
5w5feJvag/ncFHpvCr/WMZwZBz236XEvl1vi1+Fm7+RzzZCbQTQNcCSe7got7VcE3x4Q3H01eU4r
DxBLHiAZ958uE4D+FDqI65tQndMGjVhBs1HxIWSOCF90qYUfMvwFiKfsY1tbr4xo7O/peqbA/0RW
p5+Hs7wqZR+IToqmfetpBUptZXh7e4H3BBqYRZVrFfUspcTJWdueG6ErTAfeJgMqDZoXQ8GGhAD5
3V00GxAmxuA1cdSYfWxAL0Xmt4AYw316r09AASLZYOP5N5LEXS+3dhvb0A6U4SkWR7rwILdjiAFd
VSPoqY/j0E6x5JVk32QBIpWn9e+ckDvvLljQ98AuvONqqxehlmklL98EuLlNPFxenJ8BFL8clQV+
wbDxhKHNbDQyI7d3CqrRba12zwyHCSeR+sCYxk3anmtQenSJtnOk8WJXE77ps6P0Inv6tYwdsUKk
Dudx41jZ+0va+9lA81TcsSXB/XVeHm+EJ08dQfDH8vL9kkMyRHlDMh4x+lDX/f213smqFh1OkJut
XNbksVlS9yLgpjAb8h9EVxyXOMqX+T2Ia/qWDTBDDYXE6jW+wDUWZc5mQNo3h/npZ1XOTIMTXNOE
7Up6YkZNaEX8XHa4D70y87La2SLbQrXBRt8eVPdJ4k5J3j61vci6uJfhdiYSyvWPTXFZPxRmzR9s
1dIwii+xX6Ie0gYMMQnuGVVoHDnrGGkMDbl8fyRlrS4el+Cg3QZHY3coMEq7ACYgoQ9IP+2JDgIk
JtQmKHGzVQedqJhUxVN0was0QnPArW6K40ePfRImJ6py/H+uobSG0CKRXMt74UP2xbTqp//o1AVc
i26BC3J9IA8GldbR8F7Fq2bcp9ChrdqNWEGrbpIrhWt70s9rD1imhfO88QX/bj7sajVzJmH2beH7
tLYu8SJ0vtO2LvrfidUZPvq6/9KAlwYHUxmFpdUqpbz9L4NE4J03ti1bKEp89Z4m23CQi6iGhmjp
D+fAnEshnKiCjqQMKM5WN1w96TYzfiCZZUTdaf35Xi78se6/k+ceHV4vcuCdDRKbx8dqZehXvZ7U
/XeDsF7jCuNMpUIAZ2XYOU1/Wbnu6Wq2ucaGKIkXkBjqj392Ez2Xys3IMT03gt4uvUlOaOmvYILe
WO8xcPyKDAT2/7Z5b+AEyQy1vR0K539Nipdhtkl8KCAHASPSNlpi6+hzu2KG7cEW7Mi+CdykGCMm
kLOnAU1PLzbZLIB8dlJ/Uet4EXHIgPlmOg1uisKgkrU95JXXH2wC2h54/0d2inM4HyB+2zXYIAFh
yfrg2NeiR5EAFGXenD/paDVH5B9sPPG6+owNJqitO8XEPX7xMqOaM3eQrDnVG9gLOz595qMb1r48
RND5gaaDSOuo1b1+UYPpcBl5g1ik+bxBNN7efgBAs9XfK4Mpcf+MQIBirQiYvuAk4FPJY7ymyi6v
U8lURTv+mSS3MHSNt5D/22f5hkK13e984mgoBgnDfVcp5erU7eueSjzX/6EzIcYxm73aHlHrq1Ef
O5KayCEEKBR/x8mHxpZF+AvXjyRAEv1RRXQSNzApMueIPiLQI7k/QsvObcXC6XsVdE1sfdT83LjW
TmbaL21C1lb4WWr+tdGhg5f/JHoo9YuYpDb+oEiOxdhBnT6upO9ptQzdB1NJEYM79QYJ893WYwer
TaIuO877CPnEY05AWTEQuuj7a2xsHdcPdOziQYmEPeXPrXNh5UO5rMvy9sC+pVEf1zHCeT4cKOUd
eEdq94NcpS6tTTkMmmzZhLo6d4xqVFJRB7dNu8ORL58m1fwNwEMuymey3HNYcd0uGi3HtmFrHKEP
atiqyPxFDzzbhTR0Rec282QQX37WF4b5ROSHzCPAu65UmraaW+zMTS7kQK9LDI0gogy0AIybx/NK
pE18/DGvRMbBwH/6474iSN/5JS3G+N1noVACe5G3yElJJIOLKJfN7tjhMJur31DPKMXflQZy94vr
b2Eko2IEgNsmpdwXNGMXshazLBIW3ii2Gq9xnBD8BCYFRB3X46pckoTLTjGQXpIBfxR2nW2yOOiu
VEBUQQvADWxy4brZKLy2xtaCWUpPiTtdY0caYraYVLon0mMsVEBbBZMzaf2ULnyDmWVRS7yD39/H
voUHO1OkkUDb/soohm++vZSysoY+/QG1Pk60SiQkL270tyb46bLzng706Rygq7N3VtUjEar9ExPk
VqE+9rI7/a5NNajRIpiby8iiZCsdxoXk0JBxlskV9N9Npae6vhZFMvnEulTlTaCZ3bT/IQbmU95u
mvo4iBlSOfhH0jaSWKmZVDsZlPm8+vN+BYmEdg60vxkhjW9c0rcb1fI3WXkC7WyujP4KWeGiWVSO
z924Vh5ggZMpz1Zmul8/rPuROAHjMaJJAcyniIHwBlNwTYkhsJewj9lT5eyBHPwWCJW6Z+2x0OEc
bpbezx1kMXFSmHw8Sd52kUoSM3PJRO+BYfytQ5MzCXHsJlhN9ILnYC0SMxWi9uI8A5xHlGrElXks
gMSulgIpmvyMRnVqW9IFPDAypk/dEDaw17+lMYvWEar5eIgVHXz4hI0Gf6dOCD2F9wPqufcVg7dI
JuMnBHFC31EHCIcPwKtTooL6mqVJek7sYdMhhUJ92esSTWxyNC9JYEIHhPa5uM2DlYJS1tvO9PB5
bSpZHnHPAAqa0q8JiT3xS+PJGAxanTJJrYlao5klI+9tFR8vTUUrinwDZrzGajnOtcQELTAkYcGf
68XBke6YeZR+b4gMg26d1Eay9Cw3TEAtwPCsMFXI7Z6vDsNHfq99xVAjiUwpm/ImAo+ff3eBwUp2
i/S6oCZ/w0okQikEKEK/YG9Rg6tix3ydTPjSNC+5GkbM3eZbcPcjPq0jd+HmzGfwytcAJodzSlRH
4kfdLt+cCyE8+1KC+VVggzUWp0bbsnQKSVl9h2CN3l5NmROwVhbrxpAb+CfZs4LTKP6p/2SUyLO4
60xfsdCLLdSlRJmfN9PpioHafOBv0s46wN3aZyZLG16CPdKYQckmr/fCwsZ/H3qiXaC/db0m4OIU
3ESMQrpt+ZwO7Q/mXDMQKSTxB87QeroIkKwvWOXb2Z8tGKkyMbgLxef8GgXEIOAWnKVlKsdt7WP4
HARGFXJq1f7El6owVYBebFCmpZZDdXjcFiWNS26wV5anoc/C3Fy/AxIQBsZQzx08A5zYkWGjLeiT
D8iBxEUgWjMQgBhqjPaxf96BxyJ/lq8PHxVZToC9WfasgDUug8QqpLUIVbx5XnZC/u/wSgnsn5UL
2Q8rZwjifSCjpIL5fj9iJNOOZhQG6y2eh2IJNKwsb4SxQGLQlpmXk+TnxSb0phBHgry6Sc6q2gH6
piyXXEDrAe+OGk/FWaPsk5m+NaYurzsVQt/rJDOcmsbO/eoPKw3qtmyc7gJ4QFd3LkIlDzADYFkF
Wc6nlYkFXph9d3V/4pefUSTTGMspvr5jDCuEqjarqNx1Q/xm+eBIKatSNQ8yREdf/v7MgpyhZiqC
N7JLFNMhnZTba/ZoahcQzIao8oY4Jwplodco01dMbVETlJsAEVKlqRxP8lm0bYv1OoBYvgbBrv28
JUedhI4+q90Xl6FsHybyEGI4a6DwGPr2mVpzk2Ct94bvVTt040OE9fMVu6s/hyoQLHc/darYx/LT
Z6+KLLG9Mxm/bzhr830QjAaLvXJWUmk/t2U/B+RjkTe+pgkwzer/avoKULbY20AYjPEnajvTnAko
yCpl/Fhtsm5zCKwATQDs5keLkAKxHmeB0u86jgaGpV5/ZKmT1X7Me06sMPvMuMle3TkCOiZFUzqA
ilY1ZUJQrBTiy1VNzszrw0tIV2u3jLpto2zUtXKQcKDKvXRbyZy+U4kZoqoD5xizXipiqW20OSJA
7R1rrmcW/6dRif3lvAwhnZZ/TLlhhZbK4FAxCzgNzi6izOjL/a89z0xdbp5NrUheZfwthhxAvZWb
z50odZPN/kZaquvKg8ouZT2vTjMad63M6NEGxvmOtCFiyq3tlkIyxBUt7fBpg1VM1ZiSJR4XaPcK
s8v7yn4Ni38hui8eJPIWpXhMeu/KEqHi1NHpUCpWePwZf8hBRL383pbOftux8x6p76uE5kbF3SYm
+Fa4BuEUoCXefhgK8IrPl0iEzpa+yZw4+jth05SZKBBn6j4fKNhSKnsDkfxE9ZmdWU2i0o/JTecW
GcCjAdohgC6UeQ+uKDi/yMsmrHBhifvB1+sSTZLH5tA9GPtDZAix9jueqlpDmjUYl8+RNQPsXXr1
qJfjdhBwbRCcs5+Y2zuXiqF8z2XJuoOZP0tMT0oswoS/o4/OkoSxdeDvjSlHkIzsex3WdqdPI+AA
0txd0qY8i9zEhCWc11EM9v81ALACoxWNUcPAW2tl/aCWe13EjVlpHX5tOG0OXj0oxNqJdXtZjeNM
WGfjKedbHcUk1JZethGQr4cvyTaoLF6B4hFocGb3HIp7hDOg2HdEMJ9a6pD6KGQs6c1/mEVjekp+
Z94TrjIdP6dHEfGIpexJMRIOPltUDraLvbWMJTpKxEZIlO1oO8AqnC4GMeo5jeM3dJKG6ncek9sm
P8w/E6NtDLXLog46+KZiajFcp16tUY9ctouVJPgmbpgc6YCoNx5ozWsJWX75IvBVnAar82fIskAW
kx63q/ctHJ1IqT3ZoIeVKxuFJMbfriOlMHqnWDk6IyWZJgy05ko0nJR3+8a2TrFRSsKp0F3duahd
pZtemvJwluXUCzeFlyYYT+oVNzVSXXUgDMvLua5W7oAzShfEP5WNYcExnlvQGGc5zXJxRAzgZH7R
xXPf7yed7Hrn/A+20oLlkAiTc5KD0ifGtSY/Y9K1ve+BZhCzTrtRbbeMGB23Mk6OqOC9heQEyxjj
5FZSrMAmAK+Y30fPaSq4ik6BskRn3+t4gRfCiG4UOBVzmPW6gI3Fz+HV1WCm+OOIkldbkFttYiWr
suSvTaI3tbuzpO4ETVT3CJ/Zorh2topAhOp/bp+8l6ZLa6MlHolbTP2oscZcnukx3oRoLJIpqlnv
/c2fDFYA8feYG+ZB4DsUhVc3mmBy4PCZDEqocza+HjBnela/1FT5CjcGLLbipw0muSbhxc3Z6Gcl
t0jjZij4UGsb1WeF3JfIlCd7M8pHkmXMPQyxon7LeDt+yerH/XWousIFHi9szkziI5hoT1GoPVS9
jDUhNINGrau7dzee42FmyiXQHT/CRwe6Z56hoOrkVsM6kax5fsK2uHdeB1D4lyhCqOBSkzpBrEhw
la067Z31RsiFoQaUPUTf9SOR2BShsksfcOaDWThB52ORiByKUsT50ifsdIvXmUHYvlD1xkq0YMOV
Nc0xFG0XaIJtCJK9q9xH0Yd/z8uS3igdFyuqIUV2AvAbLeDuPxJeAZvRX0fXrmjttamviHxswaCT
RK4w5TFtTPgh0mvYeqtY6RDJ0QLZ5vy+MT6RdpExjEsewCYwcbElw605A187BSGVIUhs2UKUZ+5S
xpFJMYznCUdxWUPRget2L9tVNdf7omqdi3TiWq56QF3S9xv7cRM+ID0oBo1juf6k4/GOXWBImyLS
oFobcExBRlYbajn9gsIRQT4uPaAuDwViRWdM79VTH/GXXghaseVGz5k0qEyB/vVi4i/ftEsNyCmI
Mv1TnH3dBfEFCPfQtMKLFi51LguJAiO3sxAh8Gh1W1Yu/ttVGQP++euJX/oaEauO6rIGAZ/NxH/z
StxLbPV0zW8a8vekbUSezQMIYv0vbt7l8va36BlLlj+Pp7dyWHGqhOOH6Z9jF/4CPHHitEpojxLS
P7WRDHWVdRvKAB87GIjrP1oh4PvK5i8oTOKi0i+fJ0EhnEbsRkeTqpADwvPYFr4+JtwP4bdrAHWR
QLGpPRAeJvmrhmLQ3xpD4p0ajnkjDRTdapJG+OHx/xOskZDzTrsWilTTZCBrQfhQbP+5osrdR9Hs
J4sGuNckmNjiNnoLU5jucWXT8FFCYlt1Kr4BkFGyedqyzr7UMBcTdGuQn1WNiSpyqfx2e/OLQ55A
xIp98WtNM57Ghw8IRZx8p3nQkoMck6ReTfRtCF501WJd0JcuiAuHkwKG9DYQWXFcnRLLQ+KJahbA
KD2o+ZlLjGHPdzRar8My21+dSJQA3E+/AoqNDic6xA7yVpLetuDr7GaJFFo5GKLbZJgUmnWLH7kw
usXYP73XrTonYG0LnbWDGbkmKoGPgMKlu6oYMKljLCX5X8TXbIzpbGydhWB4thPxH1wCeHV7ot9S
5H/svZGMRw0rrAnGOv9tP1BZ/yIHdydNH8XpG45eC+7d1zwU7Gg7nlS7tmHMNIin35nRjR+CKQKX
PRGnHKDoXzu43vEAUtOmwlMD8t5z21CDy1MrnbUMWM2PudtP7+JQMmO0Dfac5kS0ppoG5HD1h+zY
py1pxPuvoKObd6CzVEFlwAWrzMf5VRSfIXcmrmhtlxnBrRuHCi3aoRkCoLew9SWF+YcG8AG99dep
dzWoSd40I/j5LYhahS02NfL8iU8AvZz52U/dnzwSSQZnQI2e2u4sYVChXuvwEZSW1PDiql/6gSmk
vL60gamF4LOsSXmW3WZ2PbqOzS4SCSGTYjH/ozzDf+/hIa0wmcdiegjM10lOxwd75Ym9xFNT0nop
U0WT4vcbqO+C3qOB++WgvGztgH4/wY76pIQsmLjy+/5A7rDy4seC5N65i1ccSTc2231Z0HSOoA8X
hWv05v5NY1oh6L0OHjiOY0r8Nzr1OtjauBp1lNWrrOvcfBG6Lj+EKEfF40I/po3tpfTxf2Dr2GvG
JbjB9x/IVeno5cgkf4DKZnDLspXcezIkkz4Oze6S01BdgJTfvIj+lYsE8tRR8OdqAVobkmdloi6B
xyitcO+3JzrvUw1MH/vK8xNeIpSvkB2KDmS9JYlzOHcckfzApXVb0GtazOc4ww5mBY2E+VYn2+X8
FTULd2XV+gXEfPMsIR/ZcvCG64FkxHxzgfBcv65Oro97y/nudOPLrcn3vixcmU68RPPCK2mGvXvc
Kdw8/IuIU2Zq2DNMHjUuMXnKptLgEKiAGF5JO7uVwEsF0DIblBX0YtWqOL5pLRTJRkL4c6FKIwW1
6r9i8gil7anOpXeQ5oaykkJw2X0EsTiwd1SKyzq4OAwH2Z+TfCTzZ4rW1wbdkmjJ0YHj5rtQXebI
wkzfLr7CoGx8KV4onKy5zJUkj/h8bW/SAePU1tCGgQhpM3weiIHGEeC6pbUNAyJ9YMHTSBY6yzVw
u5saQNmIyNcDE/tUNvXTooKc/vm7gwBVRpUxxRj1bkITnakC3J+sx3FDHcvNFNE1sqIwSZCmhJkl
sQj7J2ssIhZwlkuDWdDS3ntEPwUMrz2EFYzn+Pf1/r27jC4sDCJUHpRscafZCaceoLXWr5MTHsNI
5gmsPCjum1aUi6ixB3FVmM3VL6i9qbBDdZ1JnKipaDvxP1JVF2nzYHVOHC1TlJhH0/olvxXdHMgz
2FDogIRmJHyefG0CRR+R9Lf665h2A0P6ju08ozX5TLYeqm1T5LPNK2/pOQ2qt7+VMC6p4JVxSeuE
QSuUaSogafqdIX/xMku9THOxyzPXLT/UEswxFT1xBB+5+Fm4ttMXp/K3uhoaQj+EGbwBAJifQsxu
xeRThe85mOMIqYLNjHG6lNt9khm9ftzJHOrjm+5uQRMKrAYq8YmqrXsyR6x+hei38EFNF78a37Ax
Pn8rYrqTACQTaWVLMHMGFQKpszPm7JobsDbDJyI93t8gZk8OIK56GCHuoaDa2V70vWy5Ac/X/AQQ
UkVqtkf0DU8LaMQnTBB44I1+jdkDloHi8svxwOGLdylWcKY7kH2UN5IBKVgRGhQ/UxcVfN1DBB2e
wLPaBSBEaI3uncQwYUNUFNObYbEHqH66MrJZ7wF3Dq5T7Lg6yloBK3rq6xTJymbllYggEqMkInX0
O3ORsGzAzQOd0FvMxOmDF8YUaT/34iE9GsZCNBASAhq1EZaWYgH2wcYQDEI5vjRO9bw4o20FdLNp
V8aZ6dxIYNF+UxzcI8QkD2Nu2zKFy3hRAhagd7DEFaMNJta7qLv07nMB9wO6xQjSh0aHktW1pJIK
/yBCmVcbfRVp7InHQc8oDl5WLqCHplJuJTY+mWZWw+TnDjVzQ/dRPGhzPJdfLua+CTZOEJiF/sp3
v/n+sgUJL6PKKwtPp2WANpuxLDLzLcf6JjU39NYhB5NmXG69l33KhvR9WfBG+YgA0XBDoLRWPmbz
opYtfXlZeglfWBlGmqa0AsBZ/JTHEQPQHUVS5b610JoWtfMYxo+TqavRkfGX+10XxudufYuGfgVs
XCxOysnmjlGVWW467/WBMJHKtnFwn7nkAg8LrIzCtZntalDYVk+8ON0zLaiTlWoEcY0JKUHJlXHN
g6iX3Glhv9nWJN9ZlRhO2guW77gwxYdFhlmgLFtR4+lRGOpO8pOOh3VtGL7jpF0yA0+M9Xfg8kGj
lVUwPwGeBMcusgKkx3rDj1uNlVo+KD/+w4cUTzOTzTYyoTv0rvq/p7NZGm1vCzC/ZMGuDtoBzlUN
UhIfDDeUrFH5kGtRa6VnSqRScdgGddm3Tnhry6mDQHML8iE/KhJqyNWVU/64YNW6oDAwnHSY92Rn
ovNSI3PSusP3hX7lnMPJalX2NdyDGcw7l+b/xjVLMssSXCmHhC2JkMyZg8u1yCtdFtDRodL4idoZ
Ca85BH1OwZBSG+bovACMnA58/JUoud7LSf8VxUL2TYBy+pbLk4vuvi3XDETQfoKNgR3e3Gl+T4UH
ZOGt/rvuqqXcCjXL752EIGT5GeFXASRLy3pVZATuRry2tmADHU47+nZChpVDeY08u+5UqO3ez8DM
LPmENIq5iWeR7P/XuXD7nKLOSKk8bX+97jUXX6fd2qLEDHgcJiZXnwhkNbf+LQSParOwnFZV25gV
V0+ir/uVSZjVk4bQeI+/GDHqZJ5s6rUxazK/WGqv6gfESH1AmXgZaQJIZL/B+dA/COHq+Nj/mwDr
03nuG0rVoPH8ojdQbx7+STXdicx+SWr5HAcfks+PzBlJ6bAo5mDOoyBOQzK0f+k5IgK/RoDme0Kj
p+TIwmWCEaunH1WXQfajhs8xkuHsHFIeeM7UxFkPbMkU7RhD5UFnrvNsrhcC3ZnLPja7r1N5WzL1
bWFpDmnsndR1nKjc8Gj8lKEPTUw2hqoqCFfkGlc3NsxyLZEcF3RjFLyXUb+6DyVJzlRkXfnMkWJI
qhz0jlpgLjWpECyk3+Fbu+L+3ZL10F0NODq+0gDsgvPC1HW+pnAMrC+gt4PIZ1ZS43GwOchFDvgn
bx2p9b1q+uU4BZSFkYPfd5TC6Q0Xy461Gt67yCfV30NzmCFO514zGjB+MXHVF00Z5c9SbZ/Nll01
cx1+v6ie5BbjFQwq4JKJ4dU9EhAeu9xFr60OIAzdrt+aWlwNmFi9X0S36EcmLw3TXZuMvI5PbTUR
jJdTfk7aXJceXl96EfJhvu9MbG5mDLt6toanG3BUzEhmyrdUP8xp9tS/CbyGPell/+me1p0CUyBp
YeWwv0coaTjePPRs67shWMxtOlWAaTeabcmEhQmDYWWM55sAKjiTG9WlYoJrGC75/cMFg2ppwUbX
PeWII9WeBfTbOhQHiMFe/aBZQxOfWixGpAAZmmarzME7q3gRCSvFGQs6BhG+AYKpYJ74Y2xf4+AY
utzc3U89eEy/NiCP9nq9tOAsKHgHBM6xu4vW985YhCSJYTUO43KSyIJ8r0CrZBlN7Id9KuYxh07o
ha5+vULtLSHOdk54W0qapi8iXd+bI2CXaoQtV4/i4GMwvuzabM82kfSJaeyJcsXB1kDc7m7ZHb12
uWH1t1rh1jCX8KzlIJw+Mtltkv5T/U6xGzghgJ/O/bARp7tfeFu+d7Rlz4bIdlumdOX0zaIqXRLx
xf8ixpofr1sEt2aCt0V+pN5JG/8HymhDAJZaKasNicXrcyu8UsR3OIn/RJQmz/tqFOBDxyqosZ/j
KeyI68wvANbhQVow9aySBYDj1eWpzILQYgR3/Xoi+aKWQ9f839DI8pyEDPwQhu5Np/onaK9ntAk+
T3L7GXhVlfetMi2fkLuivCZykfQxeyXg007E7CuctQ73Iaj07v9gT5dFGtq6WrMwGvwYMHSOsx2R
9XUCZfIm3nTnj9JZihR9K5Gt5pNefYgtOd8jLKPbIVmyZEmRn/TvtMaxLT1r59Ao+yzv1LArNtf6
5JlSx9f53srvrJotRRtOlBW3mjw+FjW7FTFHMJeCLYhtBBDdcpDdfVCM2/KngDNxnVMLO9j130NG
ViOzpWfqqRsfBKj0XOG58DWC9AsDddC7pNbpNTeEe6ba1jE9u8LFrWBcktxD+UJ7Gls2yI8F1GSi
RxTTnjrhEbL+lkHz7aJ7vZ2HGyD6c2hHAaj9uUrsZBR9E1qZsxsKq6DKoi8DvC3pO0e7Z5S/e8KH
oxpTLdajFuZy/OVa9jx8nzZQykv48unZNWBElu//Pt95EsKlBWr5Swoe/KYnRoCHDQA+m57tq5hj
q2YA+geV+07DpUO6IzM5axXHiAc/pBrgdA9nIxkOFjh7jWPsuLHGDLwrEGeqgpPI+Wyb0C9RSlUd
L/EQ+1R+i7S9G9RV+TkhKsoHtvREwJE4oWMMdhERJHsGOg9aRcaPOw1mnBM5yRx5VMh2wM1VMpdv
6fL0wUhxD0bVLDlGR5yxQQPAswmrt09akJEjU4FbBCIlX86cRmN5FvAJT59/yNSVGiG977VFltcj
Xj/gznGkY1vfrXGzsNnxK5nnmb8iHSSv1G+SGQnO5/4dfpNPtzOTOqVxMcm3DDcqhJLK4bUILjmR
VOAixtFBOpTxTftn9fc17Fl+hk78TXtaQLIcA7PHs5YCsEJjXBDafW7JMZKMU3skvK8Hf5TpDILb
8IACSB1wivtgURadoXdMEw5wfMtF3ZIlxKnnzPcobKgJq9jFBEwo1QCG7qNdFIICiz1a1rlYoSNy
AvyoV7ii3mKo86wNn34173r2+dGt43Y42byPljSJTuZKJrVN1BkROV9wTEDcZ8+wsa3ugUn1ohfi
gZEai3OZchnXxQ/9QNorUF1pcVkBkeTXjx+Wx9POZgsCCg9QIvscifKj97wf/9HnsjeEHszNB7js
xyKODMCrRKPjQJAELUwjtoQ3KiwRmvx90d6awLydKUIvJLGh7c/CLlWqm+zu6acsOKNaPOi1Pq2l
RVrtnBRY2FbLEMVhcdXZWRHuEDd/vjqgfS5Eoboht/S9Prr6ntrKo00T1owvE/H4H9YQBaTltf0U
rx1WfwSVtO78dMOrixXXN4QzX/hYtW0OSVZft1YBiemoZqmCJo75vD2MNAR9aXfuTwzPPNma7Kat
pxOeIdwQF8qn7sAQjohTR3PBarhg4otaGHqVtIehkMNFS7Yk+bM/Njz1z/L5zw37o0GUn72CezKt
rkj6z0JQRxt07/UzwxwKHYoX88fKxMDX3UdvZ4g4AWgrI4xfFipbAkKSGqbWB3wv3WLg4Dzl1pG7
zoo4A2TBa0w5RE/BjkEnjhTZuugiOix5DsHbW3n8n/kQztgu0GQTMg1MjT4s9/411HgQEW+kpG12
A9ST5/35SezfiruDEo108Ojkbbd0eN3zXaK+oOGZgSlxCtftpYpZuO0gjAqJyyZBFz7rWUUXKGWU
2QFtQEBFZgBXFyZYNBRgULj21cDv9G6pzpVrS6TiemTrd/4rplNmc9Dx08uAVLesahsvDXMur+m9
h/axwy9CMlNmUjViljXpA+jYnZwce2+A5rrydMhztNkBa2xhGDqr95wMLMaYVPD8bdsbXEQHwlA4
1rxTrSGcjlyusSvG5vhghNddwV2qPqbwPFqe0hXxSG5Nll2UyrH7f93YC67qVPMbEfgJg4+Mx2gN
NSeSlR5Rlw4x5YWNG23mgk5hzPIYEo2QoJ5YiDR6PzApL1dwkt0YvmTuDSnrZR8Oxb35GlDphu8E
jX5T+7kk/tH2vym47I98DChd7oO2u+Zw1IXP3Ls0K7MaJpHJh7VwSIg2CWlkGHXYmYVvoqhliB2i
wEJ0LZULHB+Fe53UhV8fPj0lFr5g0IoKF95426HEFrhj9PSLS0Om7Unz37NFF+2qVfbt0h1GfdIA
94gwImGGhUi0gtTMKnk9MEWRJGUxs6pChiGfB7RfxQa7gTOwFtHx/xOe0xhBuia9uYzd6/3rqeB5
vPhGbPyr3hffvZLhhejsLrgx0aeV01GDkzZoa6XY28aDr9u/2DOACsPFvyjDB7zPGKJfJ0hIqdHY
TkmYdeKYGhOqdnjTE3CP5evJK002mMTMq+5BEX58G5duKbtzVc1Zcj0VEFP+xNAdTpdjYme1RTrM
7+JqrvzJi7Eo+TjIAq7EI7NDmENCWZ5sy7lpNc3OP29mHEI5t3ZHOUPEEzBGvTknmfDrMq/IpzSZ
mrbkcxiHTEVwbynbN9kJzUV1KPnmvg36yjgwanMOkX67pMdeiDFxO20IzrDpNlGP1wv+2sCkRcGk
bgLabgQcoTRA8EcEYEMZaCBLvmaRwe5uVlNpkik7MSHJ45pyBuXhjhwIegsQ15t8pHvlsW+kgTOr
5z8NA+a0ChDg5YhLcyweVNlImEm/JxQIaFRz6SH3DlB8CdAk2xYCsSeUv0FMxseA19fLqi0o/bgY
8meW0LUGYnuKnCNIScoGA5kJip6+JtDJkbPpDb/BCU+3V9aCEWuFmUUVy4B8Inb9NPpD/C66GNKZ
UOlY3aQthfgXPzfby8GP+lWwllbBHkIwItLNVvB0K6ynEi68pFGTEIT0RLB/ErDbryQPSkHG8ZXv
gseKlBEQmSoJMjgzBH6qAvceRtgiaaRfUfrHS23q1B9KGXF5tHvhajVHhzGx2WVWgHkTOk1c599W
rBvQLw50gh+dfkPLUDE61JrFZ4R4Cfv15on13/tMtWTH4dNEIxZRj4ykqCmY5WyrS7i2gnE+mSqQ
TTSNW4KGxbPFrUN23gyfy+0zMt4j0mGPir2zPk1aUKsktPTKn9RKFM1eZfHb7C+tiyjnpwCDzRNn
vyjDoUvxd1c5NdKCt9KzAZT+lotn5D7DMEEyPH0DZ9uN/DsGCM6Y56U/5bF2eCBy5p6WcT2/OgXM
paxmloCUHFFDvPiJR7TO+PCAQe27QcAmIS6lbifZNX0pQvynJUOpIWTupsVB+2OnJGrd4Tv6iANr
Xq2Qy4r/VIEknjAj+Ke/x1/hO2lcnkQmsJNbJx2MZw7U3jtPJxcbL9sbVjRFIzFrWTfeyIeLzcQQ
s4p+gt6pgix31usg2FXtZV3xrY+YHBdfJbZ9cdJBIkv+fFChtZTy8W1pUbut6omEOwx7lN8AnmfJ
jSeWfvI2S+1kP6vZcJi0lUvI3y9WLZlT4JTaRErbhWfbsGIVl9qPb1m+/xkws9ZXQoUUhp+ou5wW
w9jguxcy4y59U0hNWOd2RX/PuS329duglOtIRqaE0ReAZhJ0bGpwNXAR0u6InB8ehrGfWMkVBFCx
uheE7PZO/IqgOlcC1ykOZ3OWsm4B4GKhbfL7nyDTl7AwD7V+Pf0XR7ZWYerOgG+MHb4QbWvQusTN
lzRekUR1tWPEQ6Do2BkBXyP7+lpl3Ch+3jaBJ+DB5XMrLaLiwPOpkfQuhvkcj28NNjigb6W9ALOY
uzHFU6RF/H7TNfNxDnDOb8R/JFXgssTYgYmQYCnFqEP8xELvCp0UmO8JGC99sLRyf59VFyTOoj6X
r7wcGpYP7U4iHGU6MsQzceOFts3pO00b7+gFWojvFmyAGojlHgj+iLK3KuYPYkH84FxAPRnUux4r
Pq9KZsvmoO5WGPAXT2FnnOBQaNZ3RI1x3XyxG2HJ6h1kYW58trbr2E4/3y4ARZpe2exOIS3bet35
S73bSIDgg7Jd8B1NZyKSzFE4YlcEVwsNmx+h2hTX2H7ZuEljnTIsBo52+vhYV2kjTft1PwFyevYK
7+9G9NLg0yWlOArQYK7IiaeG/vgFHQhpiKv20Sl0HX+Ls5WAuzDNQfaikxOC+ocObfzRuXeMtrZn
igm2K77hrPZkK6teBK406ltQmaPMSZEwzCEmXS9fKa6iBUVzfad68IpjmwVLB4ClTTtdet6DilFm
roT95M5jlYbXxG2uZJozCWwDrpxArrzEtnQ4MZm2J4lmiFWEnB+6LrGP2WUs8g93DsQZI5T8szpH
UKZ5Xcc1CjB9YWo03l7d5ru0FDHjmd7UY7DNyvobPl4mkkbnaaE/ePk91uNHXTAaeTa4+W/N9yK7
YlDMsbVde+5l6OaiMEU8Z0mIBfPiYrCYfRcBi7foGGVtvjmcokzvCwQu5ARLX/UQr3U2eyODerch
ErHgr6dpfX9KRd141PcvqMqhVCoLzWXJ9qJUzEJa4fVhVb0bQa3Vvs0583WYVGKNPMnNoDjJgCEx
c5pkSfvlPA3isZtfuri74o3XDE4cpdignpx5BGjCtDJp+fvT1ty6zyXJXDYXdydfz5i7cTlJvzGo
kdfj8V0nOeblx9VVtUTE122ja9tZu6GcnSMAmRT2bGCAzunBMzJGEyBiekndFnhzhMvvj99ZNtmW
J1RSo5Yj68yQW2x8+zmBvHlEG7c0UtQU+ZBG+Ns3WnHfVTfXMzlD/vKe6YlhRp2agXQR/GVMhl3p
XV3nvqPYnUSVo3448F4hynsn0AAu1EK4rPD7z8HBMNnXjC1f7XvkmI+98d2J/M1foAbi7Rh4v+6N
M82q6DdT9ugaLKjZ6Ab4fyPrk2cp2HBLxTII9dwDjReCU8s0ZCm6nPBf7SVe8zamlfWcNSx5xJaV
gSEPE3/OpOzWhfEzutVks9ftuTyKvsY07gLFwmnbaqZ98huxwSS0x12ED033R0cn7tT4QEOKX5B3
toYPqfQoOjx7w9b5cjOXZlP1VpuUv2ah51kxiu8iOX4aox+KReDO2S2Qiu/7f7w5Ymi7osZ+1z/Z
+ARXSHfqIHCqJYrJZUXt5Y2I11x7uGnIkuLJTHjmfWxO0Dqxx+f8tWbp7fmuP5bl+LttBiIQ55SB
AFTk6ipQ8H3zhXO/oLJGcKv7PB8Ogzqvc5xaaySo6w+D37aWe3GKjM7JzlwrwBMcjCw1t9KDPFRG
0L3Y3wrUMi1L5h2AXaz57JNNtS+wcFwS3hnEAn6QX0cfjDl9EqPfVSr53ibEh+p3GqEA0iuSI7YW
ojCWLmsCkAcsEvfQvHUhpLaRpyjuAw/baiFfN7aASJP8QdIar8Fz0vSZLaBqd9mpsYnJcMFJocrk
8AiwlC/Ohg5AQiDMod8QS1CvXefJ7yCqnQcup9BJ3HmTHDyoavm8qdvqnlCWQ7UV228M3ZPWetjH
hTmT/lB/SxzRH/Ig27HMrpWT86+ZOohd+cZyr89NGAOAqXc0e2r1iDE56z+SAlq+bLrEIwJNeESO
c+5/4SV7GmhguM8C3pcVfle2N8HCMrSUW1kNIUXRpmXLockpuxvTHRUIWlIp0sEsQ3hqbNmk2H1W
ekFS3YNonzkWW5UdW9PmB/jevJELMUFXjRkm4IEm5WY7yMWlwfwnFmLzEVHzuv28QvIvrqcv4nwS
JBIoiwfm04A9r0iSUpv2B/kBbvqQ9zy2JUPw4DGUYH8uKPZEGsxUijQLPJlJI8Z131CVF5JuDq4g
M+FWNZyx9McO+FD7m8fos0+6Ka7jclOczSB2OSgZmkqL2P2Gtzx/ZFpIPBAWnXpG4GkAjDErP5Hr
RlVscvHZwWzWXhIEGogJzzh5wn7xGwnnro1YebCQhqHcGJGiT2xr79sen1kLJZ8HCnH8+pWTgrGW
OPr693hytTkpbNK7m6Lz9+XP0rI4HRBFiNckucJjMpyAh3xRkma6mXlljY1/X/H2bTcgxvx8ar3d
cWTdF9OiQ6/5IfgwawCwv6yqeTCgwuwhNmzQkiUBuFhw9ix9ezv0RXvz+yc5VQTS8oWxmJj91hQD
6RCaTGK+E6FoCgIAH5KZAR/5WBOQTzA1VuNKIRijvIV4v8Dpc1yGd4e+4EzJzx336N/XQP7blIEp
wH40nAKhCObottF1ZruV38bkZTBSu+Kccg1T7i0c2yh+pSJL7FwbwODYUtUwdtByXjPt6vkUhr6H
GHuekk2U7euQV1Aw93kThiiqT1q9ciIjey0JJLRwM+VjTvtZouf3YKOxLsA93GM00vqxZpXd/j1M
EtcPGfPSfMBjy+/iqfXLMYP8GzBDObOm2JZz45wRWRY2sZ54sk/ea7SU0SfH4iZO8KVHNyIAx4c8
epmoR7priDIToWRc4aK4fSdckADj1ZKiP79wgqmwBuOBxiq6kh0PwsnFAWfk1WUvfX+LJ0RrnwAz
rrAkZQfFIswub9QianwKld84bu9gFqjKUTOAIIWFChUxaIG4pdIxHMH6MnDeZ+EZgFb/OajaNDZW
vlLkGkT9XRzqU2X31DWjCfU+HpImPto7ufYqP2NnJgKNKll0xls15i69CYEMlFxOR1XhF041EVjs
FqIEhemUBloldV7gr03xRVdHmgaNz16fq4cj743j8R/zbD3mmika5C7vh9CpYeR7PWdxsUtW+v0b
Ujj1jaMtuMaOeyOQpcVkqRT7PCyV8fkzRif08HWm7OCo957CE5sjJz3j9QizWYHdsIJT6YcapJPw
xlLKrug7TcDvxJwKJujp+GC2yTbZ4OBiVcjLRZXlqhQhiI1z1jF117p2SqmmJ337ySWveKtJqfuW
/KIVzbvmHlSredPiuBqSOX/E5QNlEVZioTN8Lx5jZTEhl7R7wxQm8ixVYVpQinufYiii2KE0+zj2
qiDSNBLMpXcebk3m6h+Zr4KE/cbZzrHqcz3HlSD5gGqfDGXkVjm7C4YGeCgvk5CvJtUukmBWK8eM
qIIKZ7rAcoFLdSgPqwhHC8utT4mBb1rAS0sokvLBLAoiByqmJW/51pE6iwHcanptFP3W4p0jAwHZ
pCJK5FsUhqrp7UoCeYdZZAASaylu1+HDzxxVdo5mU/jO+eG6jW3l9LBr5V4MH9W70xa6qqZ7EhGD
GXlpvoSWvbM/uSaorDC+JwJVO06OlhR8wu3nUEnWxMq5KCTkYZrMYyQxJg468VoyDLQPVOkbW4Op
SjD8Dqcc/EMoBT4osT9o/RTgCDRiCq1pJENX0pO2AQwQmLwN/C7yx8DQ1J/1pqdxjRrZnmuUOgTA
a6FP3qqkw7PQbFD2PhDgz6KCsbz02jKCaVObRpGJyiQWHP+/iFpQtEQsM1fGz0yv2o0TYZFcOHCZ
gtoEuC+eEukWKzBVFGWk6lXW8ysMnAzd5bl9oPvfGVPXHcVDRGYYAg7TUeSvJbcsYoDGumM4A5fd
D/EMtFClda8uZw6ZfAfm4bWEef2yOHvmBvbpEGrmImGl1R0sC6oCKcoHEBYf6Fnif16sOpVOoz1a
eCnQTRsyTohGMHmKoGdUEshrXpmg2KoDX+63tqNPjRmaV+y7SpofWSty+6hNypqDHuq58yEt6hkr
R5xwmvltJVZmx+J7Qn/6qtk99aT+vU5mFNucYyNE+lNNiKNzW9h7+Y+EIFqJ1+nhgNWcYqLObVu7
0LJZvHinGcgtuXwuB+ffY85yH4YlWddz2AgGSHoR+iPssio7Xr6yF1VKTEGAzwZFw/ENyQgN1p1F
bpN65CCUuK+3DWh7oTEz2b5PtVY1DLgC8//q8nBW1hks+bbzeSqgeyMaustQCAQdvba7Af/jnRgH
MLkF2DFnjThqAi93ddcq5Qxx7CEKOV3IlVamupcERa5m/Z8dx4C2uBKFQRcMJNqvcfvTVd+0fsu/
hgrNm1aQhxjmkqTx/KKVo/iY0StNkqkLYTpE9mgxeCokZU3TnOuNYq4QSpqdnQ74qz5Bm+0V92G+
wi/9hhERLXjytwFNtAE/Yem/SlQUgCQUlKQg9QLMY1U3y63q/I1UTiAOnP9WROIe6HcyhnUAHAmd
95pWxdElmSHRUlevzzXkzPcljsL5byd3IL8WSlxoI7NeC563bldC7f1qbhR0BLNNQrah++xMakNS
wUqTtGU8SFA/6zG4v+PEJDlDsX2TjiVZ/crLAx+Qf/rgLJTAju68xUoBTCzNyb0Gqj8Se4/nqRQE
T+34oMPUNbhxB+ME1Lmmk9p6RirCzFvBT3djGePgg967okY70/vBF6O2jEJ26AkMdrKeoyS7sP5G
qtBFJl01GmWRxxMTUqAhZCzBtMZM0Hvm3/dZhcbRabLDKOEwdh/hZX+bG77/ZIywwu16kq6EGjsT
FgooiuPjdUQKtwTSvl8oCFTBKIgPGw4ubunQGn4C20rC9GXH2IU3cZH2QPOFEIPINq34vcePzGlM
gVTOG9u3KrAU0F4ibC1S5/HCVd9ZeehpMKkGFMLcfK6vrG45ZTRJiH5dDrkiewUzMkqwO30nbHNq
Eg9UAFj7IqFNjOmOJvxYIahtPOgYJHK6rgi/m3QPYqmLoVeC6e1X6z1cTuX+/RXnNwlU3DGg4Y1A
WfsT514/hDXPQggL5On0LKAcW0I5Nq6ALYkI5R8OvFM9zbkfTdbwG2bBN88EqJ5R8lb2vNKIclFx
sopCvRMCgOeqYyzwluzziMfTrOeeSP6G6PazJsXETptxFkA42Fj8hjFRusfuz6b4LiPGbwS+7Pf4
Da71P+YjQKwB330XjDkcLt1YQCGDFzfCq7jaUkcSdQ9ZnQc7zaRnYdMTADQksYbecdSUhQfRESer
kU4wgl9BV/n265w+XlVyZXALwAKWjKxGY7AnwzFpcwjIL9DFsjQb0N8IyffBWpZ96L8LSfA+BVrE
U/SNdbyQAqhx+TYn90/rWHXwXC7nxXXi06xHdFAqVLPXx1ca6TpsgerA050G2403L3Xpqk6T8FFc
fYMz1EM4f+wAGOA//629XPm4OQfsxabkM+xsFOgRm0M3c7hDJNdEOcgn4dRPMSMeqauaFog//3kR
RYu7iEoerptReiaCt3oX2Aldedd9GFOX9PfbyiFXfv9hTmwDHh72Dcsc3gLYUBbSc4q1QYLS5G3x
DZN0DANNZd0m/XsC0JN65rD8M2XpElh4LtNjVMs6yq/pRxPOm7Q6YSG++do6UPhlzPLqClpXjf+Z
vhy9npiik5OCMfunBBnn77cgxUUSm/KS2xK62VyAKbHJpOj5wuJmtnIqboC0C44IZz9qWX9Ojuly
F+YI4tOM5X4jbZYajVm3G8v8sMrC+qKYHRjQjlvDLGK/t7pKnbrScbiBTRmzxDSFuJ75msG1JcR0
i3MnCm+r34a2KZy3SCPvAAEQ8r2FTS0iyr8zvnsxggRNGbL9iooHKdrlChnH+vl2xD9CPhhDweip
K3cIAaJjbktxll4onghe+v788KZsid93PapW42ioDWknxyajqBJym50SMEkPWdoRIFTOQpgjg7SF
Z64bu3CgzYN6G7G/wGrKZsFZR5pZdOj03VxX69PGqwYcE/V+LGUVi6uTGHUDJ/2njsz8Y9ZNhDCH
3mAmOOxRHOAtHtu7qOpjxhP5GvZkd7gRio+fWYM+rhTDmDvwJorsWAih8U5+HSzVeQetrr35T+VT
CSfDfWr6wNTC1BslyXU/3EIQOrB4BnNmAQiZPHEv0rXQ4pUbdSgBr6bM9LH+LrEdVQrMJUJTCS+0
m02FmILPOlna7ncHOwWemGICDZh+dqDID1Vox7/lJpc5xZGhyiwLa1OYTBRrIT7tGZ5yLx7jf9ep
mPAALzyrEYCuMriseYHUDi1QZ8+GyUUQDCXW3qCEUzRb+cUwRtfUes3yvvlmzppxGx/1vZyVW3pk
3crwb2UnSsZQd15deUS51bX+ZJZKMWvLpP9Mf1sjdjB91OI4HxDlrpzyF+p5TqskkgBkKmQf7ai6
lcMXcKk7zwKtb1G3M/M4qmRoeMXcE1GER6gNi5tNxerPB3Gt2wZh9Xtm2uC/dPt6GqyEqM0qXtEM
avviNU+G/d/LkC5uep92jGQSbS3FUCQqWRl4mV/k35Ux87RnoxHqgWNjVBmpObZTaPeeSm+M9kER
2Z73o9EEq3kyacJB6CsTaa202F1/zDciPlBzWfXI7Tg3ekJl0JglLilc3O4OBCpfVDEHqMRoUlv2
8ZVhV2L2oi8AD8BAHNYEY0Eion3k1grgk6nqzLXETgnLNUNoJu1vdPqdA9IowDY5AGlJUdq7ER6M
iyvs7SlEhhRazxpKDY5gZ7OJfVNh2roFBRkErk3DGxO1DTJ0+hbo2GMW8kU3/N4BAV4bS8L/EcEf
e903DHzyTt2CzWwyh1a5zgvyK+HLCq3AbfmN9X9FMsE+ep6bTccFnPfySSC444sk/1B6N8Vmx6vg
P+djdRjqzOm/txxXJz8zNcJKYRYHC37YBJIjm8cAQLiWQRILIjCNRclc7NK4yg1fucyYwCWGBkmc
bejo3aX9D5eTT7EyGXcsHhO/nIQpsqejbbI2Np+Y5vTKxnbYGPgA7W6vYYw4nt3DaEW8Wr6nT9mi
DY9Bh6IjPq7PBzdk2TLwrRKVXJ2k2MaBEj8mZ76pK+sy0kkMQKgOnHwKawv+EYlbZ6fwXyvEsByy
n84w8k6QAHhf92IkpSKksRWSUOzknDaRBMYZLWxA6ODejgVq1dbrs/qn51rqBYOOrJ9RpbxVZmSM
Ht0aB+mIfu38zUvhKt5VymawxMNYout2GuukrpnBnH7//ImQP42uLy+WZu6PXdKMWvwHBFzacm0T
E2eUPE/xhs6cZKZ70MYerDuNHzniVFffvuFEFgH9Fkq/RIEjNQJn5aVRrDfksaQ+wEHewli3GusM
rFDmL2mcWTyaPKNevCfUZeVjS1X0F52+//y8gz29kjosGkF9iEBIFAUqjovedMyByjSUp+el9ETi
TJtUHFop+tClyhMQunruIJSdb3VWNb+TLoHfYhOX67NajJiYEj5GyIAk1WimyOSw8x3u6fzrM76G
wON6NH71V1+7gJafcVkKJ8/GyCl3FebTaehR4nP7mtROOzQpJ2+klG2binUFf7t1DnUG5IpsMzT/
3V5DAi8dVCj/NgX+YwLZVNV+dlfNPrJPYgP43rNK+TA5q0bq7eF50wfDw5QxIg/3o9Ua9O1Dx4pO
H5s8ZOItmXu8Osdgesfm6nrjDy20fF8bWj1fA0yUmgssnsDuJnEiiYEs7MPurgK8AfhV8mBgv/3Y
uCUF2/iue0PtB39K+YWSUNb48F7Y/2GbrobZrOXDTgSxkXfsmf0uZgB+Zj6rNQ6IlJ3cBEcCpWKd
DSYDttkRgskIfvGlgxS+/N/bVCzIcywXA2FR8eFYnhRPFJxU2VULh9t5jsM8Px4WcZ/T6xUwHVSR
U5FgHkJRXkUPXLaWR8e8R3EGLMIYPKtGQgPLdScr/6bxUr6aPQwtHyi2qwlQlVI1INSyxWOabfO6
02OPRl9Aa55wJr6NnBx7LQPgwFbUsX1MWcdoMokgzk48vSNQKGtZcdAcA+Gpu243jjwebX2EJafe
nxD1CMBH8kd3oNhsRR7fJZK1embPLhbPfQRngi+p24TrAVjbqpOuJ0WCog1NtGn5CMEPmKwtYv81
Fl1vrkuB/D2d77DaxOAY+7jybkObAWVO6kZzOG2FVJOr/uHVbWQtNxzppKjwtp3aRX4SGvmXdOxz
J3AEH1cyhwjdsp72uvIBasiCBLWog3jmXCg/A+0MR0o6dJnnUlmwEQ/ddRJlFtDWJwWm3IeJsYNy
AytFEp/2cJ4Pn7rRayTLak6brS39r77Q71XPrlOjPbflf0L/1O6cPW1cDBPcTclJBxbxLZerkViW
o5dOIRz+/4XZcETEW0/KuvCUlYVFO2FsFCHnuSmcZfOm9Dq+u9Dhyfqwg3Q5HKX03/1EjNxvWlux
KnB8TCQJgK2mDydRpp2hXWC0NxOjy6HYTHmqraOsKJhbBmC9g2OmSEBNCS5HsD0S6UCIUMG70mz/
Vk6o+50S2jy9+7swW0mSAVXjLAaoUhYwmZr0T9wg2gSs3wK3qidcGEdaNyXJvBQSpsuu2+xPE/oB
8B13n2hGIwnvgNLTV3AxJbXAIzhXSKF8gs48M+C/bjxIk7B/Dv5bgIpf8L6Dongb8Fh+b+sH/qyc
LcggzeNswZxyWZddeEGC/WEDom88YVjGtZfLEXRLiLt3B5DNrRNHn1SGcY/8E1Bi+IOmk5/s9hZZ
fmWaEaYBX2jGJagBW09z37teLQru0AxuZq8LsVa9IMqChqUKzWBIrB6lnNN1d5UGyZQcImk37/ri
4DDA97uNaSoFLjSVWla9DaPiSbObFkXIRKf+8ynECkicFQWq8tZzgv8+YtGFt5X351VO0LpS7qy/
tZQZ4QdJPhTPa4rGtCaaixGohLfwOrySwO9RmnB0jleOH7Bbh93pT7VrH8fc0EsKw5fCAEnsZuvw
/iJFNVIfpfKLJTybDkbeyXCtWkS7510XY6rJFSwERBZGLhxAbKKHl2pc4c4KTU9PG62HcTNTOaFj
2tCpv4mqaMOs2+MloxnoAzlFWUiIlTWYXjo7+Xcv36CNfPt3OtczsOePFU6YXPYr9tOcESDoQwhw
dyap/WEULToar/Gh9NOuGunnQID0zpz1qYaFxmWi9sbtwYakhM93oRNpBxARVz/xb0nh8nmnIR1O
5l56ZgFRqJyHavWupf5e+d190rfGd5ZGDfnX1RPx8W7BVSXvH08z+0c59bCDr2eCy2KlKVQYdado
E8YGs81QkR7HZ//cxkygtfc4B5M1gbcwuFu5jAG+Yg1q+YLldowl7EagVVNRGSqRCTatHfbZWs1w
kIDCfZPECUC7p22eRJqLqxEin9GQezSn0EdKl5FurBkju09b/yCmAlEB1yVcz7L0xEmSV963wYHL
5Md19nJHpJkRqwcW/kkeKlnkrpcbo/CRuFPjdK+U/7Rxm/Eh91RFsHD5C0pa62gdGCt7QFK/1vPE
VokWho1zwKJ1G/B94u/KtBupel+brczkD6PRJZzRkIFB6Y3hKarWMcac03JAwdH/ikWrgEt0WQSb
7wzC4rzBkWk/u+fQjS2Ts4lKtOnFuPDU1h7hzR2ycmUMUups1wihXz5WGU+QT2gZdSlo2zfIZKwa
UmGXzoiuCWNksuNhDARDr9NokxYOjgrxZJxIK378CgvMm1KfdQlMtBg4+t8HwJDsyMFsMUQCABcB
vcBVp9OxEE3OO/zlm0AmORccDevQ30KUcL1Z6q/Az1pdF/2x0X/dFbHCtr626dDIMhcBN083LrxJ
1fYurv9ZgIA8ap994o1aCApjG3UPaOursfpv+7lEQon7HHIcnmbxZ+3yCpy5XeAli61ZGu0i+uIY
bfGV5gOX/6aRIW6rbumlNDTtFRGYv7cDfrKKINWhbhoAiVxxRReOsVTisR3pAoO6Glz7bKFniU4I
14BnZoD6rO1sFQXtTV0EY6HWITZO4VZSC9uyPyWFaqoLgx3m2iUQsjpthgqkrMTMKa5o2kh3v6ol
sFE6lOocHPfN40E41Ri3L56uRwxeDK6Fwdc92Zhs3lWi+2rLfpwAfNskgEyBzdPjj0nfkCQxyZgn
UBFkRTbt7x2XoV+w3qYs6He7AsncaVEc7YIZURlop4GKchc5rE8enx+GflNFNjQ/yo6p4VDBO7JE
MghHqHGkmWZzH8S3M9OGkuj566hxORq2M4bpBlmZN2CQBCYtjheFnO9X+r9lJJOtVoV49Cx+HAZS
NASvp5UNm7EnPCNjysGzHcUK0amC1yp3O1pQE1s8bB9t7VIHEXEaJmxyEUCdVbsE3VA49jO2UA6y
sV9YPkGiqMUvzn+8Nft+hzwDmU7Sk1APTJ9+Dhx7eyZizmWYQfSVwfRsMiE/gb4t6N4R8npWUL+F
0k0JZJu30XCI1bDpfYgBt1NREzslwEN4N13ugUQ8zHcFWIVbYKwxwd2oaSZjyZAgXg7xbJ3gwXNY
XAXDknkxVeT1PuaFsqM2dbwTuj7ZITtaEcGKgfFVqadwr4dEUajJTsfWsJVbC1BaH+mRjN5b/21W
kdrCJHHT4lSjoJ4C9cljTo3Vctm65zwGIXT40kRTBPMF2DLDPINvAp6ndV2ltaCao+U3TIaO4wDN
2k3evZ9U9Zh5ZNPiFQ1jCCEuFGuKya6YBFu58afzUy6GNB49rx0uqt1uqtAZlsqft338xzhwz1D7
6c9NICgmKHCVZN5G1bOD6y9Hbj81Yt31U4i3FRwFNgvcayG79VxJH8EjZCBvEe5DTMbuAQv88kAF
6cIb4pVMcqtYSLZieWbEgZo7EdX6Ue6WR3fHRHMsamxiZiqIAM7x0ltOehyBz83ueIUmDkiRisWv
A7ub3vVZtDcHIpM8w4brGw66K3Fjyputqy+pM6Lu8kDCoIZuF+F4tYDs1iOGEbkdf75pol5oqDRq
8/IgVegi90j5NcHlmKuDLZB/nOnBdKFU0zBCYRkKua2tQqmKeCgyFR2gGhB3h5YpE6OnHSE7mLD6
jJXOZ4fxutAiv8DYRijhk66+46wCcxDLKfin8z5BhcEmonMKeKRh6CpuH7QslJmrCo8cgtXlz2qD
StnVeKxNxwqHKFdFoJrcAuXZtQfsgvBXaqI0/E5hirCNLl0DoO+a2Zg/ligHiHbgK4+BlgAcMISD
X56V+m+HZl0XHzNVRmP1SRoZvEQd/VsHbLmccsS8euAn1SkTi7SEippAF2HzLazs7jSmH85orR3E
C6TmcXsAE8rE4v41hygdOqSnlTsv04WgfVgaWeFNZaNNoONye2vz8MhhBWKEWfJZ/fqXAV827eaY
FyNC2zjw3TZ3CBNzSan9uQVvgkM/9awNjwrO8dOrDaWPbJb2VQdupZee+2rbci4aVtOvnO1rnhLK
yp0uwererCYKa8fS60LrGVC/vA22AnbRkmml9/O0x/T+VJtdlPqfk+FqXbUf/XDuWpGikSRii3gf
Bi4HZ+uTLcwjNmptKP2GjWSiV3PpGbAn4dhnr68PiEqMs4fDnWFEw8imebKbpUwdrlm5G4v1CrJR
0N4bXXMN4iD+NGVIy2OO42yFWlc6NaNJw3DeIOkIUREMSc1kuHLkUFaZ2YplUqt7ykE0+/35ldH0
zaRY8mW5OKwfbJMIBRRuODBEglYRe4BuYMQwagIyTczu/mtJzZCZQnYygiK29vDaYXztrg80KgiT
H4tUSMtr6tan8VznqtKaqdVlawSVbw3O6t2KIwZc3ImI3DTbcZyguZJ4N/U8nqVLJ924Fp1c0RK5
OeiKQYnLY9UU7DIdSqgpVybB3dkQOqoHg+xskMOatygNVrfzf2JfVm7+6B/3GYQt37bt2jRh/1Xv
iyvi1rhSri28nIEJzdoPG530F7kVgQGJ1Ronxe00uYqtndj2GohOnQ09VhF/ja6u294hVHg04m46
yAF1VUXjVKHuSfqWjfuMUF9IQv7Tmfauzv7w2zG+rgOYDa1UGlyVJf7VnOC7Xppvv4dG9T0aJN1j
bZdqY/XhRmypTam1vnyRkCz5S8bBGAXmkmZ4SmuHhcndJkRFcbeJlWFrDBgNuP3fYc7lheC73Okm
MyGgV7R8U95zMmYMEONRJ7IjZr4FWGn8l0GLpyvP0pvRDxiypve/MraVwCi2F+MyVOhtxHkShcuf
O5HNSLb9IX8iHEfNdDqGXgWHlNZ7xMYyFKWRt+l3Q63nlDQJAn4+oRTZ4jV1s7ATAihM0fveetn4
UnNd0BI+g5D0TGArfdO7MrJrLBq0sVZthBOqEY0Imd9cJPkM9uyF0DnGo1oyiLNKnA6HWWarKuJn
bHMuchKtkE9SQ81IUdfM4uhnrOR1zxF9laLdn0HyEzNjpUoGoUp1Qn1pGTJbqh8DkAmkVJJbjwoX
73Z8xOpc3VIj6zvWbVLisujZSEtMbW1xNuMiCFhjJ7o4005NtNTxXlW3p5f7ErqpfXx5XUkgCaFP
VBQPZnLvgcbYhWZ7WDhiSaC98QN4TRSZvO6mH2bkCUVFOJF5vdKdtWAm0BJ8r8sxvu5UvYM0Jroa
kyVS97SBrTZT35/9C7sGykmEAm7/9SAsTXPmrZSX3R+ZKO28Cx/Mn+jPheBbjb5UjSO0lTXPR5+5
AYdxDbbzL0qXk7NdF9XVL9R4N1Z2TfiSnMCbp7xLSnGqDD+abSUVEglU49pdOz1pvu7mAJRQgelJ
STeGVTUt/Eu73U18Lb/sOhAFCdNj6dflRuEd8K5oYuE0idYhHcgXeMLTRnFnb0DJTBUPRagtRZtB
DeWs7A6zIAKuwCdgvPAXueTytTwBww/11KWwjlfO9IzPMT4T1KF+Y4++tZ4H7Ce/oK8gODE0TfBS
ScjVoUA9Zk9Uc00SLMKOuEYNJiu6eDPLjI+gq95V2AmPiY3djokMWnEdsjb/k7B3jWLYw3zkHAop
8/3fHXvHj4fJ7Y+1gT7ZtfbvuRi+gZm+0g9OrV5Uw8saAUyQApm9r7MhzdZyrOnqoAD2BEq+AEqW
/vWvdUER/QuH5o7stWWaGlsObbjSc8BLh4qWuB8meSnnlM8KbRMtHXXenxavNWNN5QAtF3lN5jhB
Cn4Ji7Ls/4qTKGewfaURNavfBLuSxRQeo6xPE2XARtl2ZYFuzdm/qcBMKna7R7mw0zDyJHApSpxE
0xDnBZ9Imuhe1F2YQoBxU18hhYjKiLXR/cqyAizY1v+3fn9o3G5jTfXd0wv1NDBeKxf+ZjhlQzCf
s/S4NmP5K6UKd70x1H9pJFhb4g7/TFo8p6qfiBZQBDNVbnKrcY0MU5Au286KmWqpdl6wi8yhI+/m
1nHq2HIGghoM/Zhekut9+mYF19J/F8swKFQEpodQfRDI4oYUjMdDye31DHK0HVm82mb5iI3w3p7i
BvzJUY+e2zZ/RRosSFhW8aWfwgG6jwbALyE+9FnHsohh+87zOeKcURXFDLSJv4ykQ9bzj+/3p1B6
+MN/uigaUaCMqzQhsPXDBCmSBIGzLfDj6iF+NE5U7SeTSv+KI5r6+7hIGncHeO8Hy3wM+MVfoGl0
5Mhzb++BKboAKZrIEAkPvlEZPhcxGATFVv5PLe0iCQS5wZAcs67lrpZGjMTbqYp+oEOdqG2xOUkD
UaRUXjQFM0SlPxffUZ7thohaqXyogsUmD1wxL/IBlq8Pgowy0yVnxQELAlRSnnJNRqHl+1vJ5SF9
aAjsz7iw93x8d0zZa9XrKbHPB2wfQuIRtGZojkM4ewJW5FE6+bpRK6h35ybkIRhxSHIiPvvFVRVi
KPShCZ9/QoABQObN5++POkqXIRgWjcmM5etiRaDG6qI9E0rtpNu0Y9mlsfr6cIJCOB6Y31wKGpyo
PB3SsGu0I/KKm0XNGCu6anTuKgUDXIpPAPGjhoY6LDa/mRwSjBLnZzPN8lwt+tJY9wS+eU8k+Vb1
IjGX8rFgZ5jsr6PV5Me9DPPWHd0+Ah25hlHm7eAx+FG2YqDqwVLDzrbjb/DphJe+GrGX0BDW59m4
19lggDzaq5TexAKFkjMssJwzJuym692tlBhusUuVvES/w6jnEVZzKc8eunzUGobOI2/myc4LsJid
WnfgsaCQTM3tYcTcMKP5m3x83emcpqdyqfU4XwwyNTkBMDCci4TNIb2UBSNx0gm5TcqyZ1ITa9EV
ISunxpgkbcMQpTLrpR8IPXvP7V8KFYYRfqDl8nqvoJ351S2QesrNCqvfeQ5nlLKAschWsN9cESAx
8raRJx5+QZrQXa2nX9EiD3y5rmBWMHeJsVSYlRZhFDwVXzCF3z6zaEHE18NUFrhp7HrPAxSkZ9XI
XCwQWobf07x/K/EHvI/3cIuNqa165Pj7Yozg9o5/cVuNnn8sXB2FJhDoEb43Vx+o5TXB/7QkkMy9
pWTm3+anrd9JVV/VBl5atVqmuwqk+nNm7GcNpIxrf8TFJnoZZSqZ8PkzkDZj8Wm2IxaFRyAIHouK
qBR1Mrb9OyOuBZe1y+LhYokzB/TNU9m6zaY3l/PRVgXCD6Zr2c9lRt6kyagDQ2qaqOzFXHi9ktXm
I9MzdqURwzrJfuoD6rtN6JGr01wIqjNYfs6V/3JHfelrSrP5Q0EmedPm9j0qcJ03uCAt2ur8DtJb
l0jcQk5IL+OJoQuaZNiWq3jmCjes7AVA9rCxelBBzMd5embpeO1tUc7humVAWjKSlFxHXYSooPHP
PbbD0ZPnxZkuaQci7j59fMEn4UNPaGYmFfurLjE9/KEXY5oxtgmc5lDn/qDkZAdJ89Z8lRVPQM4L
oW8W5s1ZiXWfWXQaGNZL1tEZ0Qg9V6JZxTF0nJzILFVP7woAyf0DC4qpD0S6e2YGCuJUignc8akr
cozarWwOWv2ibc3jj2usMMjn+Cv0otr20RakgQzbeQ+NgA2K3g48+gEJZ/uFELMt19+5GJDSOYKr
SGfhABvKaHf0CL1bM7DWRkVbIA1acVs0vj/0+14VO4cWIUzUq2Iyi3YQCGYuvqN0iVdIWL6sGqkv
krMZDfvji85wppeBZNxZMTF47G9cs5Hr+l1FCkUvLBDB8PkJoDiG4aCf/y1PqI9hUHPSaEQA3qp1
lvYRr/V+aT3iwyPw5KD00xeOgDlFnhX83/SXH/RqIPLwcw2Vw/5ODqnwSwyffbHwEO/ZJf7NF/py
q0/MEmjDSOO1eAgXLMQezTDIWTG4EqH+lsLJrqE9Zf9zS5TMXvE5Z0UXDt+sjeHP/bOeIfh3HZaV
33EranHN+hjiBtn7RJDWa3diJYTslucsciRnpcUaKWLslSq8P4xHrsiXphGGFeoslw2kU+g4+ttU
01PwMJcZh5rbuZlnLB6l/gWYINwF8313+VqA440beF3R4C+vcjSBPXA41bkWJPRN3u2f1Sw5Jiyz
CRxTPHVZn7pLWw8wcPh7BlJGOFcu2bpr89ZaGg3+Js0DiLE2j1JGkXj+b0KwXnxvX8PDE0xCqQko
w9OtbnEtCLk6hqYVR9bkt50taBY+iva71HOgFCMysdEDbbDw6pTazFHBM7jQtRrFpGqzyzepHL0D
XsOGtp3JNDDdtv5RNnvOwPfrmWAFTgy6ym0ctQyHyvKsIUL7s71pzyD27BeNoRNQ3ktzL+C6QjQX
5u1YFWsJ0eJoYnW9Y7pZSCteT2hzCscGJx4bfMyl9uyR1l3FTFQCd/Ztde2MPprRnRv2rEROZm4q
yBE5CR5Q4QTu+ld8f2XcNUEr/p6t6c5/UXgiGqnI/k5/XF4RuwQcidzSOr8XPgcBh5X6eKImy/EQ
aYIi21uvFt2Vbct6++hIMJQFL6YbwZANid1ucGLT8fPonWSyOxYncxJBdszb0h9r32w/H7ysZX0Z
9SL8QA19v0tZQUIhCbw44MYg4dToZY+EIFcjpcPvZE2KbMaZr4PfQoIx87tM0VnUvW+08Sk3hM/Q
puPLDKWNEhLs07DlJGukoihwl525GrlsRa2nEWLp1mPkX42F1hYoV58F5dmDMSigN8DnGg/j2sgE
qa4c9q3eHhDusgpOmhps01K9uFAo/GtCy37aQN3iYzTxMmgoclaASgCGG7KR70QM0cjFsEmNojkE
hEZxdTl76PXIMpWma5BYeHAiJcYsKXBDr+81dDgzP+9grm1ei1GRkQkbQxY+eaKEYlvIw4UEmc/o
erE1WMYxwm6+ATSY2rCawpe+gC2zsbl1M0wxdaJIp+wPxezLl//J2nR5DpQ7DsW66cCADmgLZWlK
mC4mE65LQ9jfoq3uNkuHzy1jsc+UmbVwQz+kvc8qNuLcnQTDi6QiBIDT0oH/RDeU0g8x1wW8vMq6
+vn8wYMnyePMGm+KkFAKheNxhoi8MB2FpaQ7YMGfNjkFFJbOtHH/LcELXvvBDgL3YU3gzA8P3n96
oLXTz6j9WoSVZCTctZgj1P9FuInuR8XAYkIFZxdm4Uvju8sIGoX269Wfacm65lAclwXfeyz1EXbC
t8yTSfl7vt8WL6e623Y61mSTSVwXt8j3FATyyKB0pFQS+hVyiC5J08fgNXjMkV9G04fqfrqCFao5
vx9RYMptq7DWzlO7eVXr0wM5/M7bFYttnIsKzYA6Ajt0WA0ZIwsctqSgZ+cXilbaAmb+II0y7M8e
NmgxKQO2I7pVb9jXxArChoLvfo4uw9JU7X6vDE7n/Cj8H4jnd/+GU4cFMM5zN5/zXqstyyYy+RxQ
q9a4OdlXkR6lAmzW/3984toLpBvGLvi11Udy0YaHroLntDZuA5s+8YxVoIlp+HXYfPt0vjB3xVk1
1vqyvRYSdsllTU0Dmvxvi1tC79hDB19sOGhJkmMIYUUwjur1Kj5IpcQSQfYMEVknACYKLktefEHu
BVfb4IPQQ9TSQ3ApXPEBsmfIGh9FMpQpE5T5kIC5FhmF0heC8npB2xCfrFWwwTDvaLhTkZ19AOdQ
kNAz3KoFAzGcsrdNCUCnGYGB6K40TFsAXXOlmA22VapdqsM7qs0Bx9IkCTboa2ciMFX/HwUTrpY6
X+E5mrCR33Rlu06T3PsXLEuayryohnrzQqNMmgr85CoRlPjU9DTo28euE6+3jKoSJN4qj4i3n0zB
b34+wRb1iYKd+GdC1oTcTHt+lw2/gWXQjNtxe/p9Dndl/HkAO2mHXkpN/xGJMLwNwYau7IueurfI
fEwodSKSXJcd4LI42TdzdNRHZRiaLxe19JaUbYSbTBmftttpKYBaqZV/yOAgRjIw5D3bSHri8//W
Dt9GQe6v1vcGnLp25S0Rqi7Sn0hPAN7wrMUq7oKHvHuGQDIQGOfnIeKC7k+JWCX4QoNqpYTeajy/
BO4guBV/agbksZ0stPFdTRWDT95MfqhbyNHbp0WVDyrSplaUi5XVHa5jaZVR9TW8LLPBKwr7r75d
fP+Oqm7QgwRaCrmrYAd4ycYPnIVrkPsR9mHPNKz2mxqVpRfTvNHQ0EqU2U7sguFYqyP6zhnOx5yU
2FIGortA1OuT/yIlFKKaGAp/lhueZ+tlxC247uqqvlbmSC+dqOdyj4Ze1VwsJcXSRMXhh64t7rsc
NBQAuzvo7ccATQpC5w9TFEt3KbgPSPgixP81LC95szqI/7BVIcQg7WotPZ9+faRiE4Jh4JwqdyOB
2MkLU5ehN3rzG1SB5+gSpAfS01lkl9w4IP/3XeOHIH7d1BMirTOa/HiGnsCpNmIWeGIjORaoKOiI
fpfIm/nDC2DG2PuyYOykdsG7qifUBEBJoNw9nQ7+XuRiW1CA/wT73zbTRCypk0Sp0kdrox7iHE4j
AOgRYwx6lJLYkdVBz1xI2auSKcMaO4ZzVgQIMqrDOXrF0jADK6taSAumw0JwAPZ+44UO1K1LTDEt
L8MuJOA28WAb9Tvf0UxI26BWyfn37MMLZQNSq/UZ1w3iqZQq2qIPz/Z4qFzxELg+wB2ckGNkCjSy
dH3otPZZoEba7Z2Vc3UK2iGBDEnuEziUtBV4+NjJAvxYCiVgObksZ6OlIysQXV8Af/AJEDlEGTgV
q8Q2pLFvGq2mkYsxCOq8/QoVsoAYwVszg1uM25P2eLV+aKn0aZCPebnGKL2mPX31rWAPZ9PSKiSt
gXKDWttsPh2HzS//7dG9Fr8v58MJb1jxKTJ3zT6PoE6RqfUUG9KA74v/ubChBbLl1L+CvIO5m6Oi
PjILCqX4+/tg9/HedkyTj3bOFDDV/MSwPPIG2WLECdYspI43thFKbPNFHbikeL0l9a2nUuIgTquh
Niy7NdreDOSe9gbk012+WQZk4AjUDmebplYVYl7AgLoCpSFaPY38qtKMqIgJ44AOGZn209G6QZ/L
YeIXw1f8aBpHSax3G4RsXLoduh1vTazUkngCEk0tW98Gp0IAGDqye6341p+adQJdUETK+Nqf0rEt
8MmzO0u+jTJCp8Yu2gysorDkrbuXgubgA6h5fkB3X/qZvi+yMTKykcooTZ3b4R6Rjuex49rjJp4v
uQBIh5bLEB0tCMUA4/zr7dKHkMsCDEfx8vlORo08tG4RrX3FDxrpN5J/sgjXcLgZGXbq+Qs4J/bq
0Q9qu88Gn6Hf2uiGKBNU6AHHhlSb0QAELg0LhdxcHxkef7BQOEJHfEFqyIV4agGmXZMZDYiUqGEY
Pxi6CP0MuAple8i7yHF3xPmqii6GokcK65KcC/m99KzHXZwUNwP2niE07qxUuW9Y3pePmKPsXMIs
uSCYtsIU6mz3KG5+hSVPZFg6KpSYURupafj724RJMBX4ILrXdHeuvf2Cjj6VuxTYxpzNMEyufRv9
0ry7rr1jp8ejYaD221GytsM9YQ/m3LiI14hUTNPhcenz7wDTh+A7ccN/JEkG5zuPpHynLiYiX6r6
3Rs24xlBzikK/aLnJG3EyKDfOsS01DMYdZpNBuxCXe0kA4kmDb17/txOjXRwzGsk3mVHWc1me/0p
89+nSa707UZ2B+aAfIoaUYpgQlcgr9J+Nxu4QXm7oCwVX4lrQfJBaS0/JrMlUoYXVl21cx1I4sPV
KZoDXc+j3GKuKHwQq7SFtoNYq3eicj+dY9kV/kQ8+TB7f/BRDydf2AamrdWAMVgM6bpV4EcTRHU5
MaCks52bgU+7Xz1kxlBY6EpuzDH6OaH8KXU7F3lPXiSyZTZoziCjWbNORo+tADU+eUUiSlJRYkEu
iuo3WuK8f6V6Cin67PUvS1CbSXEEdYSBqCMMinWtCPVFADeh24O/7sC6d7lSNerR255itP09QBot
GclYLM8qZsSHaRZBBPA1EjtfyS0aaPBeqKaNt1C/qC41wTzl5pwTl7TFjj4VBzGmmLC4En/GaHLX
4wW4RhXDlMLxK14ScMCuN4NjMr8PrYxYQVXszpY76PcgBOqGcJL4HjBLsVUNY2EzRF8X1tZ48ghj
rFcovj785pZl6F3lXkHiXwFjj99K4xrGsznQxrw7H9zNAnYSHKlAhVC6w6zn0oWHwBfTqwovVQBy
AFUj61wqOSmoEvlIQ9++LnmbXp/IIkguWAtSTQ0Q+Twubp5Keso2upR2bdFVRt9/f2MqLO090coP
bVb8SotWyZrZvR49aaqyEuBGPoMSaycwBSLYsmGfFhtUzQ5zWKzL9daakKSyL2t32NPcteJI+32F
W4TDWQIl35vFecitfEERcKWaw0glu/NM/wvppqP29bEmw7mgbi9mI19kpoEYeZ4o7SlBykv5oxtS
6QcW2vHK5HtN0nwcWYF5hFOdvujpamiPhFsV+WNhqLLVoybuohv1ZVTzgSkI1VkGt5UFDq32SSTC
PZS8hivkZ/cIPXU3pGzb5jhMzL1GxU9cgw7mGlifuOmq+dm4rfEGefsdrdq8qQVAfD2LxFswHuEF
ioKatKGALBLxosG1vVTgH+A3y8HS8C0PDHWde0DXyhzFiuVMS+h7CsP7UMO259onwK5GqOyhj1B7
n507kNO3t6iOxg724nXwaafpYKVwnOPs+wN/XrQ3q5JQ7oGE7sZuRq0R+Uo+ssNcR1hP4PbpHxgE
gIvQB0WsFgKIPKBUzbaBYb/e/vG1aRTczJPuo0lnaC0ffD+sh1DH8KghajamXHCO88lDf+yIEe1Q
lQxvizQ84Nc5AGhXwpsBNgUZI75b3w+T2jn5Q1NDToEEhjFE2SInv+u/W/c5fbes7gHT8IzLaLxO
yn1dYD1/LFAjSc2oNdA9yy5+dGGGbKG9k/phdsgBXoiFVTLskuZndXN1KXjGd64Q2RvyFOWn1nRw
jM8VwLPGW0FbngkgaLo1k7LDX+LG4qQ8etxM2XVPeaCWdFcX9pHzM54659kLc3ifKGH1uXfM6kHy
k8spgZMqovZvVExOVfHUYvUDawcDWTh7X0bPtrvW4Uw+r4uP0lM0VF4bFRfNyHFrH05Aw3e25ZYB
NPIpQzp14GMorRb//m1EmWLysmfudgQ8+pVf8w1rPfmVbofNVkM5T/ZCVWL8zch8PK141mmnyPCf
6LdEYf0qwrTIT1hPZyg6igw/Dl2OD6xgL7JUcUX5RzV38xfYCb3ZYBmm1ovU7eZtzMrVcy4y+OgO
ebNjY60h2zt5rmAOC696f1bsp/Zg09CFlNUkU2BLcm33EZ4WUM1LWeISjDHPtJw1qnzp7EnCh7uz
u+z4nM0T42QFzTI9u5luWy6+f3YGXnoXeDt3MdLnA4dEayQiikBlrSiLsmTPvm+eWK0V74dRtevb
SG7J7IQdmxJGL0Mk3ho0AY0Uwv+0458k5f2/dlVZIJLUjDwxMvcyy+PFhEHPfCKhVCtcQHrHW5VW
Tbroc04zbVR3Eciiql5H1/6/aby1Mr9/iC86ejvI17bpKODRvsW4683XKs8U7kadmx+DA3zTOGV/
2CSpmhnuiuXUZvaGPTmp7tWhkSsyh4FcZVIc2f5HRCa+pz/7nyC6Uw4Us6FPVV+gRuKvkIuQ3FN3
qrmJInhh24YgiHZOnGeEQILGo0nMVTiDOAsKrfo/Avga59TGEW9tH97mZD57qLk5qQPLNEbwauAS
PRvIBNJYZSonGsY3QW7xN0762lEVLFWmcF0lTcDPADVQSfyA/S+O2iJc/yK2AXYv5zh2EBjzaVA7
LWosY6j76YOGS02E7hm+FBXozn/QJ1LrKM4IKG8TSv3jTQ2yBPrZGT8eUSn1nSdetCbpybZKdCFC
NztWukebKSoukjypUk0lShGxVsPoIyEkiKizQ3fN1X1JTmfd9zLy0chqw8vqaeX4tO1p7xHIycdV
ZVItvcMKLn0iT0nUODPfnlbl0V2LU9blwM2SD4CSc/Olu4ELrfPqLOOJii1rw80OTggrCf65BnLM
BNiwX1UKh6wZjnVPsvvWaVT8hifWC0KFhzVAeq4wzLhH80kUfoD06/lVhfiPU2v0R4Szp6MLx7Ls
r662SA7/wWmsXl9WBlfgIDO7p0lgfn2wmk+wfeNqX2diBLAk8n+sJY8L/+CCG+H0so46/Ic7zVGL
+63+xiSO16T7H3d9eVcVojCvnoXVVW4Af0SfQLuILqjB3bA7tGTAyG/3ZDUMf639HyWtTv0TXRmh
wiYFoJOhmnQ7WTeGPbYRO76EDf5MK7csKNQl7SkaDRbPoIkYP7+Xy0MymtROyb/n1dAPQJET45Ir
tdidUIZv9Ju5GgyXTNlgOoGtzLIHXa1kYWGn29zzXAlXMDOnpZRQj136GLtkI5HCsWmd5iiYTBX9
TNsBMXKZxCJAzS3M9f5lZTm2b67CgqF82LqtpebimubZhboOyFepl+JmNAWC7lBBQvoYiGhd4jZy
hYmOYY1uQTwvcwotpn5Fh9Bhdf463m1v29XnGhjnxT0qUS0RATp5T24lJSwM/V1pnCTPmuGG5AVO
dFfcGg8TARh9g701WBrJs6GYaN1Dg13eKs2Oogvm2SfGsJ/gCuo1ugtwU/ZXj5sT5OlX8wxpwlDv
tdI3+/Zdn06ITn3QNzuChixtdYq7ZosH5+zRCiTMzJdYeHeAn1PtZEm+s8n+sMHzay/wh8yOVCyl
1k9WVgWcoSoC+FnV5MLC2x7sdIBZZX8DJZ/0AsHZ9mfda2hfTtMHiXQoqLQHqVoSOoCcRUMSKAHW
aKVM34yxSlpBJ+hJgGXFCpBNIN8L150N9cXbXumRTOJZKxnf83j4UBmCBrRfMKgZPEdkehVSDb+9
Z/gV50XHvif8Mo29+MrOpcIPvgxOYXGV6DzfMRax6mTsfSG3AAaNm9UhU+eIQDFImCU1Jg8aDv3W
vzFk3d7W6cuv0/CpC/TCKDl27j9bTY1i5CG9kfgYKWPhhRoYPeJCdcXYgJ14k2c8sWQQZRk1az6/
gVxlSXzjwlAj5M3W/3Gya98/riGka1+qYJhv+TTIVAxKfTX0D6Hq0FWJ7ZI4L7w2mDzjTj6WouZB
Fa1h0iT25hT3dgpxcpvMhnMqGUtn9CsZ/tkHbhMt4dMJ1HJYLxr21WNmDsZ0VPXsOIoQtWeLlKJ6
63SvFmJeAJxXC5GdUvnxwXMzrL5Ixg27Wj3EO+0M52yfIlfJTuz3K8FXbxqPe0GIK53zaos4gxut
70sllhUVlxCtFu+Zko2WlJXPtcGXhJgfYtRgKV6uibNskiioEfAZ2BRhgIxr2PWAvKpnjO0o1xg0
cf7mtxe/BpY5X1MegT0kxBgfsOgb6teJ4oWNduSTLpekvG0morfsNMi4S6+uC3gSyp8ffNwaKljJ
TV+e+wXnLeM3hCJXpjxH1vZqsAb636lrhGNH0qDEyBDslM+kIowMv94kciVORONm//GbjZXlU/91
4YyzfYPahoKXgdXacy6gsRFF5CzUH1MSgsFNmcPyuz09EZSMqpXtKOhBM2jHNWaBNgTnbAdttpPY
1ZX+AJKboFAGEKHHG5vTeVpe8jk5vPjHBGcK3WO+sTfvcLYVt3PRoSTDMnqY+EwB+NJxZX+/Ftes
aCLosQOOVT+v4/gHfRldH+xhl8PqYZABCqr6hz4n/l5QS6u2tH8Nd1f7KMUO93tgl9zjiASjjtBj
soZD3jialQHcT/PrZIS5ftKfhcxSsGd2QiYVi63QfMRdOW6CmNlqDmz5XWSD+G8wQJJzCPi0baYJ
31ZsCBrqvRx4b0Xs9RvlGcUZUNmD95RsgUrgbtk5Jhfe2RFJBeLRmatvR6a1W8pUMUtxfzUNJxKc
cI7jyL5uBIVGwgaKY/LQHl8tlnt3AOYTi36/kQjEXfAiK1et+WA3Tt1cEQByT+2GzPuXrvI0ok8+
YONkphz53hYOZVYvdWxEXYiDzYzkR0OWcug4RvWHey3twFbmIv7vI8K9Fzl0ZgnQ0NdfwQqt7yS+
M3P7qwtfBJ89fnv6sb9R7PuUGHwPpRSIqmBu8EowSszVcvdVVq1vFBLmXKQAPoPn7HPBqS3MMDI9
VuK8NottAkHK1fvABCri72B85JzxCPp7pUL3x8jB0TvHyg3Aa/zOPcxTvjJGx4aZvCOR7V5A48rX
OYZ9AlIGrxexT17oQcHOtsEB4PIM/qB8qSVBzMoWo0GBEfxEIUwnFWg42yvdw4jNurc0ryJdEy49
hf3q+hkRHpNLzpyp26ecnsrPvO8QSQyUKlo5lNI1X0gCn/LhWSohTG3wdFHTAJO7dJMMRzqrkWI2
1O1OO9d2RN0zFdm0P48/SCHgKlvVsiELjHpU18YwPZFIxqyxPQt3uHdJfYnIEPNX8ZouV3ynhhSh
2/UK9cYMCZpxkWLCF5WJSQS6v4eYgTJKPXLl9uJs7y4ePgz+OfdMSd4iYZqYWhoqeImZJyes02XV
bMiopVdv1Wd75DmNJfVjtZEKIG8VNoox0benXj/HCMdI/oN2kWXan8W4hLYEk9SfoF/ESd4NqwDl
8jW14D04iPIdy/NZriWSdOC9484fTDRUnPzgMM84xZjxY4uA3Ladxv6KxxlLbfDl3xXV3gN9kuWo
r0NyKUY6WgeqPWSw7j4NeDLTQZWQ0TbbIup7bVzjK2jywSTFqCL7gDNmfKQhTF+1zvEWFR8jECqS
HrZQ9lH4b9SLczL6i9EoraWl67GrKStZo68+adk7u6D7VzgQ9NCtAr4PWfJRKqo9zZM1ITpE1Cz/
1hmebI0un2AFyFsH0gI7/DiVvz4aD+thdbCPUfRZvTkGp2f+IRGYfpaZ5A4Xnqb+7zFfpPRJM55T
UVbt9JbCDN0NMPCzHN+V+c2pQ38P50M+F1GTImNJzXMLcn2IpgvM0ZBop9Ae9AuOoPOk3CfK/ChW
UlfKZ3mlk8y2ZezqoKe0WPiKRQIwFDKPoHhCuKigXzprg1b6m8wCM8JRbBAuVVCln+wRmgMMb3vZ
+sAL1n8cOe4CdJrsZl+vn3KPvVdn1teiHREy7D1/+nz/esnT6PckB9ID4aOu0Ebd4xpNrqPnvtZX
PSH6WtC/HnZBuDtMz/ZZB7qQnalEZ0vEAHEdBi8KxpO/Kg1cs4cj0TUqOZX74ObFsj82LhEfNpyY
S1+Xk4zZaeXf/AIT6ySlQgrnOUBMEZ5jZ6RpyLld0JQy+Lt0w7dTaFz0BO4S3TrKY7gVR9kgErd3
1CuHvCz7kQ0TgCxS+rkorDJgbIfKNaUz5BESpV8EnL7sKGNYTxb0WwKrnmxud/tl2R/nvznRkCyu
Htf9dz/zVjRYEBZoWPKweCcxaLWEZuQtFLr0aJSnrCYyCswYBVVH/GNiBooj+6ZRN6crs7kg1gBQ
xqYQKnAvEinT/Ir95yuTEH5spS3bN2Q/A2G9mkyWW4RFX20PYWoUCLWGyFskBcEbMGPiFkJ2nprY
+qF8DdOtOERHm29qXqepzKZeJpWn1VdVQSGi95IzJBm693oSS688ulybW42Q9FNuyFYzwWN4hkrE
W/f6g8i5+G9Y0h8YTNPrRUdIUOIkuqyWDglQoCaCqvbGXhrQdU1SWnmG4N/xhLCL+R0ZwGiHXHHo
GfgxsqKGiy5xfr/X3qbgCDez2W2Ln/Pmc4jCtl4raaOTUDlubp5KMUupoYAQz7cNjtF9NrkGh7ig
C559unPVRFj5VUqLC2x3xPK/MByjOk1KrZH4Se8tWhl+SwbP1/v+wewldPxul2pvuFT+j472JP4F
GuP8VMXEIQNE3r3IVasuns64gwmI+t8Rc9F23ePdJjPzvJbKDeTwA1OfJP0WJOPOhX03ACptP57V
xaYTQ5wjvbtLEyZumqtcFqmhbUIgAMu6uWYwQZofuSumtLxwvhjzx1rR0FV7T/XmzsL9zl0mcDK3
NLnBCGmfA9tpLzb1wvkPeKSd8Jj2CKQHl6WKa0n0u+2fCG4ynN/fQyrT2Mb9pRk0qOSFf53wxMxL
FFNpb5A5m+kvXvuk+ewSaz06x1S8loalU7vV/DArLUrUJrtMtOqdbOKN8/mSCX1EkgngCxMcEGo7
okMxNb4iZ8ac9GHsHJG3tWogtZieGn3HxuCDrUclMNFdzBHlQPqKSNkicYiXy5sDnn/I8Zv+wUFB
2QFGv8xvOL8T8e/rX4cy5PkkUh2ptlqejv8hfroVa5Y9QUSwyNKAR0+97ebQR02xpDs/7XqMpVc7
aejzjgDzLlBjakiibUOHE3sGsZc1dGlyE8b7ZVmPIDSC0m4DiFUvb0BWlAhc3n5E7x4yAPsfOX+h
YD8i2N0DQbrhIJbDXr701peedAzrOgl2kJ0kqo/kEyoi/v59g/Sanmh/n81wed0/wnD06XQ/VBNs
eoqI9lLebeOY5wYoo4datFlqJkftOEHP/28awaTSYxTMzMZl9MngRjn5WUkc2+ibOICVuQkgwLXq
AQEBKN5FZ6HA+WLEIWvvZOS5LjUDgRymrlOS7hCtdHn9U4D3BevN5Wnsnm3OVrufRCiTsjgNew+x
LQFTHbLRw0IDtQC3my+PrjWaf2UX9HhUAjdbabVymIl2htROMFcv0ReZdGt11LUECouJL44KmH3m
FI9dyCfOQSDn4Ba8SpKSaj/VzGY288Y8/gst4+jFVpT4OLgQgrko8bu9fWGS8KCKGAPRopyS/uxM
0V6rQiZAFO06j2SMILNnVqn2BD5qHqORri8A2xK34RFbATjWB6wD0Aj3ESt26LZWOdITTwKB01sV
p+6ymDuT2m3kJtK6bxghcptljaMqQFErNEvqVns/RPL8Qc1ITiz1U7te3CS+7NOB0AtPAEmdrZfS
acSNaxXVPraFDYhm8+nmlOpz0wG8ncPIzwEaIrHr270maq0aOfgDFpyG1vq1RS9El6/XosWmZHvW
nDFLY5l0Rbgloe9XCPgjXCShQ0jAbJOqxf4JMH5shWx9YPj4R5Gy5SU1ANz6mwm73LeILDCGXs9b
xTNr3TM+vLu8Y+CemJUw2iSh8FrzRF0n5DZR2WGUZNDItTrcZVPghwvguTRoUZuf8PgRhCl9tuIt
OoHwIWffoGNBC9/N04f9y/KaCyWcAa9o/whaDRDA8mvb2Oq0/+43msHvfhjfeewvzmSiP23dMg56
tp+nrZZWmAsaBt0ZiXdz7FHcpHsp9V1FphgRIPNG2ut/MFTR98m9Hcp3XWaNtne8vXaLVqq0nXTZ
vvqPX3Kxz+bmZrqcYly8PPLB5S07uGWW706//W+2ZI874dmj1wKIZVm8U8Hns7iW9oNlEruoN94B
abXJVhj3wuwLej7yJRecuWXaSJMq3dDwXMIxcHCvkGwkNi+Zt/Ah6TjNiLhA03cJi/sSFFyoDKAS
jvfcXhL5N+uhupiROBkrnQMk8vrVoXGne0oCod1m1hZGOSN/SAC2mBQji5gB0NQ3TWuD60hgYych
QZiyRn5EsFFaIsEc9Mimz6mSqUyjG7xhuh99q9sp59ZRmXZ4BMzY+eb0Pg12DVLO/H7bYRwlSo6N
tdSPbD9n75SSuVZLnetbg0ENYzqZQnhHEdFgIJjexO9yhlvtVBsLLtVFJhOUmqfzQ9FbMgowGni/
QZqZD0Gw8NMidmzq3JNRZamtxyrLpdnhwKhvbJNBNQ24vPlVZZ0O1d2Pxn6K4Yk3OhTNU165P7I+
1zLnjmuDDZqmC29j3x/PuzEILcsmttztAedWA5qHxZJNP35Bv5iLRqu4bDBYOuNnCr5zBwKO+F6a
/i5PFI4KmndkcjGb1Qfx7HCfCPl0Q2ps1HUrWRBTiiJwmguS6qQemk+60mAl/0mbx3Aeh8FgqT/c
Wf6RP9hTrOH9RzBmBv3pp9K+bLzIzODsSXzRHGwnL8itarXZxVU/2RG7qn3NBqAJxrReQUjeJ8I/
B9uUzdV+RDXspN72mchUaljhj6gdRvqbqFvjAcmm4MUVCLWeizSqQIml900GIFslGD1EU2aUgqQt
h1CpNNyB6zb2i/IZIb7MTghGpPgYRZD24Yi53Byuzo4zMWNvSPga7qeH5U+fgDyZFWoyWXK1YpEh
0oemkjTOS4/0ajARQhJgnxSrbYXQ/VOeLyde8U8iDfGw3URVhmJo+hovX+e+x41uAX6RTJTSUHte
QxxGm1g5tgEGhelkXKDdhy21NblKtjRDU8htbv3hUdKo+9eSLuxXQjqHi+dH3g0NoMv0itvkiMYM
tkO8XPbW337vi48kJcE1KFolaS85dnTMIj3oeBBCs88EFqO6+aDqoBvgjLATbetctr+Rw1MEYRkq
c+7+731khptHlHhwv0WhIQd8Gq3Lv3ummIpeaBQUE9dNKniS2buP90kgX7YbGwaMfPDLCUfs1Ler
GtuS842DlhRTbHH46oplev4XyU3Z1Ulyv8RQD2DxV80h8de1EoNT2wKLjxeTYa/2snqX5GBuJHjv
8CeCX4b6zJkwi3wCIvAgJE4pDEqxTUi8gAMt/t9cmBWr1MgoW4lAlwye0bcHl54XIwkhF6M07OKj
8WeNmHYGsD+2KuxfbmBOBpwlG2dOSJMqwOpj1wGHGUXh7/xUAzoBo42VvLd519kTYNmPZRAElRVA
L7qrdVVyKYHRKAptlqJiJpE7T+C9BEua62M50M8bFPdTI8cDhTTH3ezfCTmQqNF47p/+ha4Jxebb
6ktNDyh4HFySQlYMixYjV9GVn+Qz6hkWlHJ8Gby+zydra2uFeieZ+x4y4H4b7v3KHF7cEnvWexIc
eQvn94otBBbKN4KYQh1bptFPjkIBwkxdTu+uRF3k+g3UCkRxyepjmKaiDx2bX7bmzP3HydQSTBlk
g7gB0han2RXnMhUpPajBb8CrGB7qb1Xjn/0BRdlblpgmH7u2EZ6B0B5ltuguVXI+NOsjUqj+93L1
RlPkMjwiUOZsM+Fa37p4KSQGwCf5vsogSJhcH8s+pismG7v1Em9jTHPTRh6Jntq2cvKfq/FO7rAM
tv4Afq+EkOdgNIYDnx4kBIZaKWG5Vc/qGa0TFzVKblK4aUm7Y2HdzZ2QixXHjysiaccIaDwmMcnx
Xm6Epz56Piiq/t8ORVCC5wYNnkhGBawiUosRkxZa0XqTWdDUUqfIVjx5F6NgmObP2J34jXce9sIi
anIimVYYDdcIkIQvbaxaIcyTneIogfcvZdsBRgrTY7MRtgIOpAc2Cqylkt1JBtcf4vOkDO+lwpzV
r+LKwVL0d1/RZ8oQd/fJnzGIgBlf6BvFzKDMPI24OvX7vT1JrAOJTft6odhXlirK30IKKB5ye2pL
1Jyk4uglAdSU3OSQkBkvEImfIlQBE1ZR7fCO6CN1G95e6GxRZGaQ+8kRTqW5w3g2hLKXa2xX4QMF
UmPzpC9jLKn3QQydaA+rKOLuO7qd4kmzYmDciUmMZwwCr7Z5Q6wiWngZ2iMCxnAUrQYEMRMQd7to
Kl77htH4KNciiuoASkdGCosXH/nHkFEfCVb+js6kYsYf2e22jvDa7LhJndCmywRTCDRhBfWH/i8V
O8sHg2z8mMQo2S3JDHYaLwa5JIH5tg7TxfKFhRToqlHT56dhkOkY6sghysKlzHCy4W7Yr/goRg2v
A3a5B9paLpEuVm22nTerRVYVeCd8uSwF6uzsJU3qWu6da4pcf86A5uHPj2flEcxm84KFMyqVaQ6A
VOXxzi+I5YIieTYYgOI0NixO7kpvBFMPxvhdtyKdcqu3gz28aqya5WCucnM8tEWaYKVNTJ+rOljo
vs2XoCvY+XqhG0L9ib8ikphjF2eieuNjkbDCWLkG7oYLgcoefCvuIH51AaADJjL1gvRMXs0SGvvS
AcNv1R5+tMXsmUUUDKGL20C+mjNpDYuG/cePgdkwZBeb+jHJoUQtkRFMW+aidwsITxqGvS7Vxc4/
It8ha0kK2z4wHAY1CtSWH9+AsEdzm+HyUZjKJIoVH6y/JwIRYSq6vOMGdWKFSO5fj2cEp1jF805Z
otUMYFe3BXqXsmy4j6iWXGa4ZITbZffc51mZDxXUloCvpyC9G5Zkhg8GED4nYzcquKpQDWOWO+U5
xJEYCXyO027BZ/paaKiasynsMPfZOarVxauYqGWA5HtEFuDsJ/gbH+wDT9D7CZ7kBDXGwwCtZrgl
UkcqfmdCTFLBU0p+Vjd8/Hh7UX4g9P00NRQD7UDqi1r8xuVcl5Md0gEu7VHD7HutghzoaMAWdlc4
MaUOk7CNHLbLhBHXdUZgS9/hxmz6hFEAZGcjqYkY2wwIDyYbbY2LqFcRbTtGPht29+OGkWU3Boii
xVc/J9r0p04y1J2dKonlwxTCgXv9XU+VwySiSM9nCAjK3eoqZiTGfiHePISBOO+k+O28ebdHelsH
gVwwXeRxNK9KcFkUtXccAwbheAULPXuSq5+g6x9qcJDpgaU6i/4H6+dtv9arDmIAf0Uh9DgeXZ+f
0iz5C9c7eii/fXDyoTEo3Gb/t8Y/EdKQA/CH+cki8F1kmlMWovnAJ/FCsENcaPXAEK+NEm47MbHf
/S0OOGZFhkTJvxEvgD41lkWy253pGiwNIsN02XKrZ23RbMjBkHq8UNBLQhuyA8uJT72AY3JOerqX
X9mx9MpmZBGbzIk07WEd7UFisk07tWDmwnkpKe1Xlknu9d8FRGLgNdXK3z8zQXtygKvqrueoC0Vy
CPOzKHJbuLvcHSxAVNRmEdORlGtnrMYZ/PG9J1N0m5hXcV5ULPnL73jOkl7/K0YX3iL6MC15Auji
b2MFTGjpMZVjoFytwv9VaLLrWsOGr87JQn9D82cvzBBPkAdP7sO1/Cs/xUQU6Zgx50btHqVIQU8v
QKBqXg6X49JoA9gH3JNFbIRG9GL4jsc8Kiz+e83dI6Y4nTeS+9HfjkQFafRwWdo9qPljeIQT3/yh
7b5IB3iQq171aHD6CGc7G91Nz4afQNw/r7akUst4sOLHFUQH5r+iFasbAV39yD8tjWMEBT2B13Wc
3YH4GlJhbMeF++d+ei1LTLE7MvlrBK98DXJ7IoecJ7GJ3WLjHGjFLQWxvDZiKw06fM61QoHRWuwF
vP9DFmRd7eIwj+eflRTh0Yjd7F92+9P2iMmOLuTuULjFXWuscSuOxW95onj8efFBDTSrAumqNK60
d6u4H0DkX5vQIA6mc0D7t7Ld0qTsN8rYffRECgEhwaJoXzEmFyxwp4n78OOIwfnyTumkt81p/Yjd
ZvqMwF4hcr1lqVGcMMUbXgATGBVU67RCdptzGHjj4xNn+ITcCmQ8v8EZUb3tc1fMJPgq77wvltDx
aHZHr5FdY3RqfGDDbED9HknmqfpEkTohkcUO6Vg0Y5PtzYeE6vI8XaCiNeEEgylx+Fpx+yV8zehP
7x9EjP6vk5cufOVZ3baALLEzOIm2GkLdOO3KVd54vT+PWwlwd19HTAQmrED4Qr2peR0RNsq6PvVf
99Gnr1ct17FkxmOFT04EglZmLVUGGtwS1xxJQyQkjMKln5Ys28OD/OCQMkJlgUQ40QDUuXyjBx89
nmu+D5JMGV2lUfh/7TRWW5zeuMT9kgzcNRAbUnL0UxhGhCW4bkGohlX7ZPVp5hr+ITuGZJeixrTy
1jk/v0aWw3I9CJSRvQLIHzawrYzKOuh8qFU/wNzIGcZdYD8nPRQAN6fbvkBXMjZpNIFSqdICxGki
dKgQAeF637XwekBPEJerVrMh+nkiHwtrUcX5MnclOn0AjKu4D8aXh/k2a8+pU7ZJ7AOY7ly6689e
64J43vSybWEk7FWi15flnwVaPTNi7Zpvkt6AaT+Y65uwGY1HBVLqTisVWRrgBHgB6k5TxuecDIdj
SQ1M4qIl7MZv1t28zRn08IS9zgN2vxGgx8YQ7zbE+HdRAgEbLEMC8JODOH/yhjMucoVewjdmDLG6
wtw=
`protect end_protected
